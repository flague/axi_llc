module axi_llc_status_reg_wrap #(
    parameter type reg_req_t = logic,
    parameter type reg_rsp_t = logic,
    parameter axi_llc_pkg::llc_cfg_t Cfg = axi_llc_pkg::llc_cfg_t'{default: '0},
    parameter int unsigned DataWidth    = 32'd128,  // Data signal width
    parameter int unsigned ByteWidth    = 32'd8,    // Width of a data byte
    parameter int unsigned NumPorts     = 32'd2,    // Number of read and write ports
    parameter int unsigned Latency      = 32'd1,    // Latency when the read data is available
    parameter              SimInit      = "none",   // Simulation initialization
    parameter bit          PrintSimCfg  = 1'b0,     // Print configuration
    localparam int unsigned NSets = 256,
    localparam int unsigned NWays = 8
) (

  input logic clk_i,
  input logic rst_ni,
  // SW interface
  input  reg_req_t reg_req_i,
  output reg_rsp_t reg_rsp_o,
  // HW interface
  input  logic [NWays-1:0] ram_req_i,
  input  logic [NWays-1:0] ram_we_i,
  input  logic [Cfg.IndexLength-1:0] ram_addr_i,
  input  logic [DataWidth-1:0] ram_wdata_i,
  output logic [NWays-1:0][DataWidth-1:0] ram_rdata_o
);

  // Internal structures
  // -------------------
  typedef struct packed {
    logic [DataWidth-1:0] tag; // Tag field
    logic qe;               // Valid bit
    logic re;              // Read enable
  } tag_reg_t;

  typedef struct packed {
    logic [DataWidth-1:0] status; // Status field
    logic qe;               // Valid bit
    logic re;              // Read enable
  } status_reg_t;

  typedef struct packed {
    tag_reg_t tag_reg;      // Tag register
    status_reg_t status_reg; // Status register
  } cache_line_t;

  // Internal signals
  // ----------------
  axi_llc_status_reg_pkg::axi_llc_status_hw2reg_t hw2reg;
  axi_llc_status_reg_pkg::axi_llc_status_reg2hw_t reg2hw;

  logic ram_hw_req; // HW request for the tag store
  // Address translator
  logic [Cfg.IndexLength-1:0] ram_index;
  logic [Cfg.IndexLength-1:0] ram_sw_index;
  logic [NWays-1:0] ram_req;
  logic [NWays-1:0] ram_sw_req;
  logic [NWays-1:0] ram_we;
  logic [NWays-1:0] ram_sw_we;


  cache_line_t [NWays-1:0][NSets-1:0] rcache_line;
  logic [DataWidth-1:0] ram_wdata;
  logic [DataWidth-1:0] ram_sw_wdata; // TODO: define correct width
  logic [NWays-1:0][DataWidth-1:0] ram_rdata; // Read data from the tag store
  // Remap hw2reg and reg2hw to the cache_table_reg_top module
  // Make the signal compatible with cache_table_reg_hw2reg of cache_table_reg_pkg (autogenerated by regtool)
  // reg2hw q and qe coming from the sw need to go to the tc_sram
  // q and qe have idx, that is the cache line. Need to translate into the ram addr

  // -------------------
  // Address translation
  // -------------------
  // Use intermediate signal to have more readable representation of set associativity

  assign rcache_line[0][0].tag_reg.tag      = reg2hw.tag_0.q;
  assign rcache_line[0][0].tag_reg.qe       = reg2hw.tag_0.qe;
  assign rcache_line[0][0].tag_reg.re       = reg2hw.tag_0.re;
  assign rcache_line[0][0].status_reg.status = reg2hw.status_0.q;//status_reg_t'(reg2hw.status_0.q);
  assign rcache_line[0][0].status_reg.qe    = reg2hw.status_0.qe;
  assign rcache_line[0][0].status_reg.re    = reg2hw.status_0.re;


  assign rcache_line[0][1].tag_reg.tag      = reg2hw.tag_1.q;
  assign rcache_line[0][1].tag_reg.qe       = reg2hw.tag_1.qe;
  assign rcache_line[0][1].tag_reg.re       = reg2hw.tag_1.re;
  assign rcache_line[0][1].status_reg.status = reg2hw.status_1.q;//status_reg_t'(reg2hw.status_1.q);
  assign rcache_line[0][1].status_reg.qe    = reg2hw.status_1.qe;
  assign rcache_line[0][1].status_reg.re    = reg2hw.status_1.re;


  assign rcache_line[0][2].tag_reg.tag      = reg2hw.tag_2.q;
  assign rcache_line[0][2].tag_reg.qe       = reg2hw.tag_2.qe;
  assign rcache_line[0][2].tag_reg.re       = reg2hw.tag_2.re;
  assign rcache_line[0][2].status_reg.status = reg2hw.status_2.q;//status_reg_t'(reg2hw.status_2.q);
  assign rcache_line[0][2].status_reg.qe    = reg2hw.status_2.qe;
  assign rcache_line[0][2].status_reg.re    = reg2hw.status_2.re;


  assign rcache_line[0][3].tag_reg.tag      = reg2hw.tag_3.q;
  assign rcache_line[0][3].tag_reg.qe       = reg2hw.tag_3.qe;
  assign rcache_line[0][3].tag_reg.re       = reg2hw.tag_3.re;
  assign rcache_line[0][3].status_reg.status = reg2hw.status_3.q;//status_reg_t'(reg2hw.status_3.q);
  assign rcache_line[0][3].status_reg.qe    = reg2hw.status_3.qe;
  assign rcache_line[0][3].status_reg.re    = reg2hw.status_3.re;


  assign rcache_line[0][4].tag_reg.tag      = reg2hw.tag_4.q;
  assign rcache_line[0][4].tag_reg.qe       = reg2hw.tag_4.qe;
  assign rcache_line[0][4].tag_reg.re       = reg2hw.tag_4.re;
  assign rcache_line[0][4].status_reg.status = reg2hw.status_4.q;//status_reg_t'(reg2hw.status_4.q);
  assign rcache_line[0][4].status_reg.qe    = reg2hw.status_4.qe;
  assign rcache_line[0][4].status_reg.re    = reg2hw.status_4.re;


  assign rcache_line[0][5].tag_reg.tag      = reg2hw.tag_5.q;
  assign rcache_line[0][5].tag_reg.qe       = reg2hw.tag_5.qe;
  assign rcache_line[0][5].tag_reg.re       = reg2hw.tag_5.re;
  assign rcache_line[0][5].status_reg.status = reg2hw.status_5.q;//status_reg_t'(reg2hw.status_5.q);
  assign rcache_line[0][5].status_reg.qe    = reg2hw.status_5.qe;
  assign rcache_line[0][5].status_reg.re    = reg2hw.status_5.re;


  assign rcache_line[0][6].tag_reg.tag      = reg2hw.tag_6.q;
  assign rcache_line[0][6].tag_reg.qe       = reg2hw.tag_6.qe;
  assign rcache_line[0][6].tag_reg.re       = reg2hw.tag_6.re;
  assign rcache_line[0][6].status_reg.status = reg2hw.status_6.q;//status_reg_t'(reg2hw.status_6.q);
  assign rcache_line[0][6].status_reg.qe    = reg2hw.status_6.qe;
  assign rcache_line[0][6].status_reg.re    = reg2hw.status_6.re;


  assign rcache_line[0][7].tag_reg.tag      = reg2hw.tag_7.q;
  assign rcache_line[0][7].tag_reg.qe       = reg2hw.tag_7.qe;
  assign rcache_line[0][7].tag_reg.re       = reg2hw.tag_7.re;
  assign rcache_line[0][7].status_reg.status = reg2hw.status_7.q;//status_reg_t'(reg2hw.status_7.q);
  assign rcache_line[0][7].status_reg.qe    = reg2hw.status_7.qe;
  assign rcache_line[0][7].status_reg.re    = reg2hw.status_7.re;


  assign rcache_line[0][8].tag_reg.tag      = reg2hw.tag_8.q;
  assign rcache_line[0][8].tag_reg.qe       = reg2hw.tag_8.qe;
  assign rcache_line[0][8].tag_reg.re       = reg2hw.tag_8.re;
  assign rcache_line[0][8].status_reg.status = reg2hw.status_8.q;//status_reg_t'(reg2hw.status_8.q);
  assign rcache_line[0][8].status_reg.qe    = reg2hw.status_8.qe;
  assign rcache_line[0][8].status_reg.re    = reg2hw.status_8.re;


  assign rcache_line[0][9].tag_reg.tag      = reg2hw.tag_9.q;
  assign rcache_line[0][9].tag_reg.qe       = reg2hw.tag_9.qe;
  assign rcache_line[0][9].tag_reg.re       = reg2hw.tag_9.re;
  assign rcache_line[0][9].status_reg.status = reg2hw.status_9.q;//status_reg_t'(reg2hw.status_9.q);
  assign rcache_line[0][9].status_reg.qe    = reg2hw.status_9.qe;
  assign rcache_line[0][9].status_reg.re    = reg2hw.status_9.re;


  assign rcache_line[0][10].tag_reg.tag      = reg2hw.tag_10.q;
  assign rcache_line[0][10].tag_reg.qe       = reg2hw.tag_10.qe;
  assign rcache_line[0][10].tag_reg.re       = reg2hw.tag_10.re;
  assign rcache_line[0][10].status_reg.status = reg2hw.status_10.q;//status_reg_t'(reg2hw.status_10.q);
  assign rcache_line[0][10].status_reg.qe    = reg2hw.status_10.qe;
  assign rcache_line[0][10].status_reg.re    = reg2hw.status_10.re;


  assign rcache_line[0][11].tag_reg.tag      = reg2hw.tag_11.q;
  assign rcache_line[0][11].tag_reg.qe       = reg2hw.tag_11.qe;
  assign rcache_line[0][11].tag_reg.re       = reg2hw.tag_11.re;
  assign rcache_line[0][11].status_reg.status = reg2hw.status_11.q;//status_reg_t'(reg2hw.status_11.q);
  assign rcache_line[0][11].status_reg.qe    = reg2hw.status_11.qe;
  assign rcache_line[0][11].status_reg.re    = reg2hw.status_11.re;


  assign rcache_line[0][12].tag_reg.tag      = reg2hw.tag_12.q;
  assign rcache_line[0][12].tag_reg.qe       = reg2hw.tag_12.qe;
  assign rcache_line[0][12].tag_reg.re       = reg2hw.tag_12.re;
  assign rcache_line[0][12].status_reg.status = reg2hw.status_12.q;//status_reg_t'(reg2hw.status_12.q);
  assign rcache_line[0][12].status_reg.qe    = reg2hw.status_12.qe;
  assign rcache_line[0][12].status_reg.re    = reg2hw.status_12.re;


  assign rcache_line[0][13].tag_reg.tag      = reg2hw.tag_13.q;
  assign rcache_line[0][13].tag_reg.qe       = reg2hw.tag_13.qe;
  assign rcache_line[0][13].tag_reg.re       = reg2hw.tag_13.re;
  assign rcache_line[0][13].status_reg.status = reg2hw.status_13.q;//status_reg_t'(reg2hw.status_13.q);
  assign rcache_line[0][13].status_reg.qe    = reg2hw.status_13.qe;
  assign rcache_line[0][13].status_reg.re    = reg2hw.status_13.re;


  assign rcache_line[0][14].tag_reg.tag      = reg2hw.tag_14.q;
  assign rcache_line[0][14].tag_reg.qe       = reg2hw.tag_14.qe;
  assign rcache_line[0][14].tag_reg.re       = reg2hw.tag_14.re;
  assign rcache_line[0][14].status_reg.status = reg2hw.status_14.q;//status_reg_t'(reg2hw.status_14.q);
  assign rcache_line[0][14].status_reg.qe    = reg2hw.status_14.qe;
  assign rcache_line[0][14].status_reg.re    = reg2hw.status_14.re;


  assign rcache_line[0][15].tag_reg.tag      = reg2hw.tag_15.q;
  assign rcache_line[0][15].tag_reg.qe       = reg2hw.tag_15.qe;
  assign rcache_line[0][15].tag_reg.re       = reg2hw.tag_15.re;
  assign rcache_line[0][15].status_reg.status = reg2hw.status_15.q;//status_reg_t'(reg2hw.status_15.q);
  assign rcache_line[0][15].status_reg.qe    = reg2hw.status_15.qe;
  assign rcache_line[0][15].status_reg.re    = reg2hw.status_15.re;


  assign rcache_line[0][16].tag_reg.tag      = reg2hw.tag_16.q;
  assign rcache_line[0][16].tag_reg.qe       = reg2hw.tag_16.qe;
  assign rcache_line[0][16].tag_reg.re       = reg2hw.tag_16.re;
  assign rcache_line[0][16].status_reg.status = reg2hw.status_16.q;//status_reg_t'(reg2hw.status_16.q);
  assign rcache_line[0][16].status_reg.qe    = reg2hw.status_16.qe;
  assign rcache_line[0][16].status_reg.re    = reg2hw.status_16.re;


  assign rcache_line[0][17].tag_reg.tag      = reg2hw.tag_17.q;
  assign rcache_line[0][17].tag_reg.qe       = reg2hw.tag_17.qe;
  assign rcache_line[0][17].tag_reg.re       = reg2hw.tag_17.re;
  assign rcache_line[0][17].status_reg.status = reg2hw.status_17.q;//status_reg_t'(reg2hw.status_17.q);
  assign rcache_line[0][17].status_reg.qe    = reg2hw.status_17.qe;
  assign rcache_line[0][17].status_reg.re    = reg2hw.status_17.re;


  assign rcache_line[0][18].tag_reg.tag      = reg2hw.tag_18.q;
  assign rcache_line[0][18].tag_reg.qe       = reg2hw.tag_18.qe;
  assign rcache_line[0][18].tag_reg.re       = reg2hw.tag_18.re;
  assign rcache_line[0][18].status_reg.status = reg2hw.status_18.q;//status_reg_t'(reg2hw.status_18.q);
  assign rcache_line[0][18].status_reg.qe    = reg2hw.status_18.qe;
  assign rcache_line[0][18].status_reg.re    = reg2hw.status_18.re;


  assign rcache_line[0][19].tag_reg.tag      = reg2hw.tag_19.q;
  assign rcache_line[0][19].tag_reg.qe       = reg2hw.tag_19.qe;
  assign rcache_line[0][19].tag_reg.re       = reg2hw.tag_19.re;
  assign rcache_line[0][19].status_reg.status = reg2hw.status_19.q;//status_reg_t'(reg2hw.status_19.q);
  assign rcache_line[0][19].status_reg.qe    = reg2hw.status_19.qe;
  assign rcache_line[0][19].status_reg.re    = reg2hw.status_19.re;


  assign rcache_line[0][20].tag_reg.tag      = reg2hw.tag_20.q;
  assign rcache_line[0][20].tag_reg.qe       = reg2hw.tag_20.qe;
  assign rcache_line[0][20].tag_reg.re       = reg2hw.tag_20.re;
  assign rcache_line[0][20].status_reg.status = reg2hw.status_20.q;//status_reg_t'(reg2hw.status_20.q);
  assign rcache_line[0][20].status_reg.qe    = reg2hw.status_20.qe;
  assign rcache_line[0][20].status_reg.re    = reg2hw.status_20.re;


  assign rcache_line[0][21].tag_reg.tag      = reg2hw.tag_21.q;
  assign rcache_line[0][21].tag_reg.qe       = reg2hw.tag_21.qe;
  assign rcache_line[0][21].tag_reg.re       = reg2hw.tag_21.re;
  assign rcache_line[0][21].status_reg.status = reg2hw.status_21.q;//status_reg_t'(reg2hw.status_21.q);
  assign rcache_line[0][21].status_reg.qe    = reg2hw.status_21.qe;
  assign rcache_line[0][21].status_reg.re    = reg2hw.status_21.re;


  assign rcache_line[0][22].tag_reg.tag      = reg2hw.tag_22.q;
  assign rcache_line[0][22].tag_reg.qe       = reg2hw.tag_22.qe;
  assign rcache_line[0][22].tag_reg.re       = reg2hw.tag_22.re;
  assign rcache_line[0][22].status_reg.status = reg2hw.status_22.q;//status_reg_t'(reg2hw.status_22.q);
  assign rcache_line[0][22].status_reg.qe    = reg2hw.status_22.qe;
  assign rcache_line[0][22].status_reg.re    = reg2hw.status_22.re;


  assign rcache_line[0][23].tag_reg.tag      = reg2hw.tag_23.q;
  assign rcache_line[0][23].tag_reg.qe       = reg2hw.tag_23.qe;
  assign rcache_line[0][23].tag_reg.re       = reg2hw.tag_23.re;
  assign rcache_line[0][23].status_reg.status = reg2hw.status_23.q;//status_reg_t'(reg2hw.status_23.q);
  assign rcache_line[0][23].status_reg.qe    = reg2hw.status_23.qe;
  assign rcache_line[0][23].status_reg.re    = reg2hw.status_23.re;


  assign rcache_line[0][24].tag_reg.tag      = reg2hw.tag_24.q;
  assign rcache_line[0][24].tag_reg.qe       = reg2hw.tag_24.qe;
  assign rcache_line[0][24].tag_reg.re       = reg2hw.tag_24.re;
  assign rcache_line[0][24].status_reg.status = reg2hw.status_24.q;//status_reg_t'(reg2hw.status_24.q);
  assign rcache_line[0][24].status_reg.qe    = reg2hw.status_24.qe;
  assign rcache_line[0][24].status_reg.re    = reg2hw.status_24.re;


  assign rcache_line[0][25].tag_reg.tag      = reg2hw.tag_25.q;
  assign rcache_line[0][25].tag_reg.qe       = reg2hw.tag_25.qe;
  assign rcache_line[0][25].tag_reg.re       = reg2hw.tag_25.re;
  assign rcache_line[0][25].status_reg.status = reg2hw.status_25.q;//status_reg_t'(reg2hw.status_25.q);
  assign rcache_line[0][25].status_reg.qe    = reg2hw.status_25.qe;
  assign rcache_line[0][25].status_reg.re    = reg2hw.status_25.re;


  assign rcache_line[0][26].tag_reg.tag      = reg2hw.tag_26.q;
  assign rcache_line[0][26].tag_reg.qe       = reg2hw.tag_26.qe;
  assign rcache_line[0][26].tag_reg.re       = reg2hw.tag_26.re;
  assign rcache_line[0][26].status_reg.status = reg2hw.status_26.q;//status_reg_t'(reg2hw.status_26.q);
  assign rcache_line[0][26].status_reg.qe    = reg2hw.status_26.qe;
  assign rcache_line[0][26].status_reg.re    = reg2hw.status_26.re;


  assign rcache_line[0][27].tag_reg.tag      = reg2hw.tag_27.q;
  assign rcache_line[0][27].tag_reg.qe       = reg2hw.tag_27.qe;
  assign rcache_line[0][27].tag_reg.re       = reg2hw.tag_27.re;
  assign rcache_line[0][27].status_reg.status = reg2hw.status_27.q;//status_reg_t'(reg2hw.status_27.q);
  assign rcache_line[0][27].status_reg.qe    = reg2hw.status_27.qe;
  assign rcache_line[0][27].status_reg.re    = reg2hw.status_27.re;


  assign rcache_line[0][28].tag_reg.tag      = reg2hw.tag_28.q;
  assign rcache_line[0][28].tag_reg.qe       = reg2hw.tag_28.qe;
  assign rcache_line[0][28].tag_reg.re       = reg2hw.tag_28.re;
  assign rcache_line[0][28].status_reg.status = reg2hw.status_28.q;//status_reg_t'(reg2hw.status_28.q);
  assign rcache_line[0][28].status_reg.qe    = reg2hw.status_28.qe;
  assign rcache_line[0][28].status_reg.re    = reg2hw.status_28.re;


  assign rcache_line[0][29].tag_reg.tag      = reg2hw.tag_29.q;
  assign rcache_line[0][29].tag_reg.qe       = reg2hw.tag_29.qe;
  assign rcache_line[0][29].tag_reg.re       = reg2hw.tag_29.re;
  assign rcache_line[0][29].status_reg.status = reg2hw.status_29.q;//status_reg_t'(reg2hw.status_29.q);
  assign rcache_line[0][29].status_reg.qe    = reg2hw.status_29.qe;
  assign rcache_line[0][29].status_reg.re    = reg2hw.status_29.re;


  assign rcache_line[0][30].tag_reg.tag      = reg2hw.tag_30.q;
  assign rcache_line[0][30].tag_reg.qe       = reg2hw.tag_30.qe;
  assign rcache_line[0][30].tag_reg.re       = reg2hw.tag_30.re;
  assign rcache_line[0][30].status_reg.status = reg2hw.status_30.q;//status_reg_t'(reg2hw.status_30.q);
  assign rcache_line[0][30].status_reg.qe    = reg2hw.status_30.qe;
  assign rcache_line[0][30].status_reg.re    = reg2hw.status_30.re;


  assign rcache_line[0][31].tag_reg.tag      = reg2hw.tag_31.q;
  assign rcache_line[0][31].tag_reg.qe       = reg2hw.tag_31.qe;
  assign rcache_line[0][31].tag_reg.re       = reg2hw.tag_31.re;
  assign rcache_line[0][31].status_reg.status = reg2hw.status_31.q;//status_reg_t'(reg2hw.status_31.q);
  assign rcache_line[0][31].status_reg.qe    = reg2hw.status_31.qe;
  assign rcache_line[0][31].status_reg.re    = reg2hw.status_31.re;


  assign rcache_line[0][32].tag_reg.tag      = reg2hw.tag_32.q;
  assign rcache_line[0][32].tag_reg.qe       = reg2hw.tag_32.qe;
  assign rcache_line[0][32].tag_reg.re       = reg2hw.tag_32.re;
  assign rcache_line[0][32].status_reg.status = reg2hw.status_32.q;//status_reg_t'(reg2hw.status_32.q);
  assign rcache_line[0][32].status_reg.qe    = reg2hw.status_32.qe;
  assign rcache_line[0][32].status_reg.re    = reg2hw.status_32.re;


  assign rcache_line[0][33].tag_reg.tag      = reg2hw.tag_33.q;
  assign rcache_line[0][33].tag_reg.qe       = reg2hw.tag_33.qe;
  assign rcache_line[0][33].tag_reg.re       = reg2hw.tag_33.re;
  assign rcache_line[0][33].status_reg.status = reg2hw.status_33.q;//status_reg_t'(reg2hw.status_33.q);
  assign rcache_line[0][33].status_reg.qe    = reg2hw.status_33.qe;
  assign rcache_line[0][33].status_reg.re    = reg2hw.status_33.re;


  assign rcache_line[0][34].tag_reg.tag      = reg2hw.tag_34.q;
  assign rcache_line[0][34].tag_reg.qe       = reg2hw.tag_34.qe;
  assign rcache_line[0][34].tag_reg.re       = reg2hw.tag_34.re;
  assign rcache_line[0][34].status_reg.status = reg2hw.status_34.q;//status_reg_t'(reg2hw.status_34.q);
  assign rcache_line[0][34].status_reg.qe    = reg2hw.status_34.qe;
  assign rcache_line[0][34].status_reg.re    = reg2hw.status_34.re;


  assign rcache_line[0][35].tag_reg.tag      = reg2hw.tag_35.q;
  assign rcache_line[0][35].tag_reg.qe       = reg2hw.tag_35.qe;
  assign rcache_line[0][35].tag_reg.re       = reg2hw.tag_35.re;
  assign rcache_line[0][35].status_reg.status = reg2hw.status_35.q;//status_reg_t'(reg2hw.status_35.q);
  assign rcache_line[0][35].status_reg.qe    = reg2hw.status_35.qe;
  assign rcache_line[0][35].status_reg.re    = reg2hw.status_35.re;


  assign rcache_line[0][36].tag_reg.tag      = reg2hw.tag_36.q;
  assign rcache_line[0][36].tag_reg.qe       = reg2hw.tag_36.qe;
  assign rcache_line[0][36].tag_reg.re       = reg2hw.tag_36.re;
  assign rcache_line[0][36].status_reg.status = reg2hw.status_36.q;//status_reg_t'(reg2hw.status_36.q);
  assign rcache_line[0][36].status_reg.qe    = reg2hw.status_36.qe;
  assign rcache_line[0][36].status_reg.re    = reg2hw.status_36.re;


  assign rcache_line[0][37].tag_reg.tag      = reg2hw.tag_37.q;
  assign rcache_line[0][37].tag_reg.qe       = reg2hw.tag_37.qe;
  assign rcache_line[0][37].tag_reg.re       = reg2hw.tag_37.re;
  assign rcache_line[0][37].status_reg.status = reg2hw.status_37.q;//status_reg_t'(reg2hw.status_37.q);
  assign rcache_line[0][37].status_reg.qe    = reg2hw.status_37.qe;
  assign rcache_line[0][37].status_reg.re    = reg2hw.status_37.re;


  assign rcache_line[0][38].tag_reg.tag      = reg2hw.tag_38.q;
  assign rcache_line[0][38].tag_reg.qe       = reg2hw.tag_38.qe;
  assign rcache_line[0][38].tag_reg.re       = reg2hw.tag_38.re;
  assign rcache_line[0][38].status_reg.status = reg2hw.status_38.q;//status_reg_t'(reg2hw.status_38.q);
  assign rcache_line[0][38].status_reg.qe    = reg2hw.status_38.qe;
  assign rcache_line[0][38].status_reg.re    = reg2hw.status_38.re;


  assign rcache_line[0][39].tag_reg.tag      = reg2hw.tag_39.q;
  assign rcache_line[0][39].tag_reg.qe       = reg2hw.tag_39.qe;
  assign rcache_line[0][39].tag_reg.re       = reg2hw.tag_39.re;
  assign rcache_line[0][39].status_reg.status = reg2hw.status_39.q;//status_reg_t'(reg2hw.status_39.q);
  assign rcache_line[0][39].status_reg.qe    = reg2hw.status_39.qe;
  assign rcache_line[0][39].status_reg.re    = reg2hw.status_39.re;


  assign rcache_line[0][40].tag_reg.tag      = reg2hw.tag_40.q;
  assign rcache_line[0][40].tag_reg.qe       = reg2hw.tag_40.qe;
  assign rcache_line[0][40].tag_reg.re       = reg2hw.tag_40.re;
  assign rcache_line[0][40].status_reg.status = reg2hw.status_40.q;//status_reg_t'(reg2hw.status_40.q);
  assign rcache_line[0][40].status_reg.qe    = reg2hw.status_40.qe;
  assign rcache_line[0][40].status_reg.re    = reg2hw.status_40.re;


  assign rcache_line[0][41].tag_reg.tag      = reg2hw.tag_41.q;
  assign rcache_line[0][41].tag_reg.qe       = reg2hw.tag_41.qe;
  assign rcache_line[0][41].tag_reg.re       = reg2hw.tag_41.re;
  assign rcache_line[0][41].status_reg.status = reg2hw.status_41.q;//status_reg_t'(reg2hw.status_41.q);
  assign rcache_line[0][41].status_reg.qe    = reg2hw.status_41.qe;
  assign rcache_line[0][41].status_reg.re    = reg2hw.status_41.re;


  assign rcache_line[0][42].tag_reg.tag      = reg2hw.tag_42.q;
  assign rcache_line[0][42].tag_reg.qe       = reg2hw.tag_42.qe;
  assign rcache_line[0][42].tag_reg.re       = reg2hw.tag_42.re;
  assign rcache_line[0][42].status_reg.status = reg2hw.status_42.q;//status_reg_t'(reg2hw.status_42.q);
  assign rcache_line[0][42].status_reg.qe    = reg2hw.status_42.qe;
  assign rcache_line[0][42].status_reg.re    = reg2hw.status_42.re;


  assign rcache_line[0][43].tag_reg.tag      = reg2hw.tag_43.q;
  assign rcache_line[0][43].tag_reg.qe       = reg2hw.tag_43.qe;
  assign rcache_line[0][43].tag_reg.re       = reg2hw.tag_43.re;
  assign rcache_line[0][43].status_reg.status = reg2hw.status_43.q;//status_reg_t'(reg2hw.status_43.q);
  assign rcache_line[0][43].status_reg.qe    = reg2hw.status_43.qe;
  assign rcache_line[0][43].status_reg.re    = reg2hw.status_43.re;


  assign rcache_line[0][44].tag_reg.tag      = reg2hw.tag_44.q;
  assign rcache_line[0][44].tag_reg.qe       = reg2hw.tag_44.qe;
  assign rcache_line[0][44].tag_reg.re       = reg2hw.tag_44.re;
  assign rcache_line[0][44].status_reg.status = reg2hw.status_44.q;//status_reg_t'(reg2hw.status_44.q);
  assign rcache_line[0][44].status_reg.qe    = reg2hw.status_44.qe;
  assign rcache_line[0][44].status_reg.re    = reg2hw.status_44.re;


  assign rcache_line[0][45].tag_reg.tag      = reg2hw.tag_45.q;
  assign rcache_line[0][45].tag_reg.qe       = reg2hw.tag_45.qe;
  assign rcache_line[0][45].tag_reg.re       = reg2hw.tag_45.re;
  assign rcache_line[0][45].status_reg.status = reg2hw.status_45.q;//status_reg_t'(reg2hw.status_45.q);
  assign rcache_line[0][45].status_reg.qe    = reg2hw.status_45.qe;
  assign rcache_line[0][45].status_reg.re    = reg2hw.status_45.re;


  assign rcache_line[0][46].tag_reg.tag      = reg2hw.tag_46.q;
  assign rcache_line[0][46].tag_reg.qe       = reg2hw.tag_46.qe;
  assign rcache_line[0][46].tag_reg.re       = reg2hw.tag_46.re;
  assign rcache_line[0][46].status_reg.status = reg2hw.status_46.q;//status_reg_t'(reg2hw.status_46.q);
  assign rcache_line[0][46].status_reg.qe    = reg2hw.status_46.qe;
  assign rcache_line[0][46].status_reg.re    = reg2hw.status_46.re;


  assign rcache_line[0][47].tag_reg.tag      = reg2hw.tag_47.q;
  assign rcache_line[0][47].tag_reg.qe       = reg2hw.tag_47.qe;
  assign rcache_line[0][47].tag_reg.re       = reg2hw.tag_47.re;
  assign rcache_line[0][47].status_reg.status = reg2hw.status_47.q;//status_reg_t'(reg2hw.status_47.q);
  assign rcache_line[0][47].status_reg.qe    = reg2hw.status_47.qe;
  assign rcache_line[0][47].status_reg.re    = reg2hw.status_47.re;


  assign rcache_line[0][48].tag_reg.tag      = reg2hw.tag_48.q;
  assign rcache_line[0][48].tag_reg.qe       = reg2hw.tag_48.qe;
  assign rcache_line[0][48].tag_reg.re       = reg2hw.tag_48.re;
  assign rcache_line[0][48].status_reg.status = reg2hw.status_48.q;//status_reg_t'(reg2hw.status_48.q);
  assign rcache_line[0][48].status_reg.qe    = reg2hw.status_48.qe;
  assign rcache_line[0][48].status_reg.re    = reg2hw.status_48.re;


  assign rcache_line[0][49].tag_reg.tag      = reg2hw.tag_49.q;
  assign rcache_line[0][49].tag_reg.qe       = reg2hw.tag_49.qe;
  assign rcache_line[0][49].tag_reg.re       = reg2hw.tag_49.re;
  assign rcache_line[0][49].status_reg.status = reg2hw.status_49.q;//status_reg_t'(reg2hw.status_49.q);
  assign rcache_line[0][49].status_reg.qe    = reg2hw.status_49.qe;
  assign rcache_line[0][49].status_reg.re    = reg2hw.status_49.re;


  assign rcache_line[0][50].tag_reg.tag      = reg2hw.tag_50.q;
  assign rcache_line[0][50].tag_reg.qe       = reg2hw.tag_50.qe;
  assign rcache_line[0][50].tag_reg.re       = reg2hw.tag_50.re;
  assign rcache_line[0][50].status_reg.status = reg2hw.status_50.q;//status_reg_t'(reg2hw.status_50.q);
  assign rcache_line[0][50].status_reg.qe    = reg2hw.status_50.qe;
  assign rcache_line[0][50].status_reg.re    = reg2hw.status_50.re;


  assign rcache_line[0][51].tag_reg.tag      = reg2hw.tag_51.q;
  assign rcache_line[0][51].tag_reg.qe       = reg2hw.tag_51.qe;
  assign rcache_line[0][51].tag_reg.re       = reg2hw.tag_51.re;
  assign rcache_line[0][51].status_reg.status = reg2hw.status_51.q;//status_reg_t'(reg2hw.status_51.q);
  assign rcache_line[0][51].status_reg.qe    = reg2hw.status_51.qe;
  assign rcache_line[0][51].status_reg.re    = reg2hw.status_51.re;


  assign rcache_line[0][52].tag_reg.tag      = reg2hw.tag_52.q;
  assign rcache_line[0][52].tag_reg.qe       = reg2hw.tag_52.qe;
  assign rcache_line[0][52].tag_reg.re       = reg2hw.tag_52.re;
  assign rcache_line[0][52].status_reg.status = reg2hw.status_52.q;//status_reg_t'(reg2hw.status_52.q);
  assign rcache_line[0][52].status_reg.qe    = reg2hw.status_52.qe;
  assign rcache_line[0][52].status_reg.re    = reg2hw.status_52.re;


  assign rcache_line[0][53].tag_reg.tag      = reg2hw.tag_53.q;
  assign rcache_line[0][53].tag_reg.qe       = reg2hw.tag_53.qe;
  assign rcache_line[0][53].tag_reg.re       = reg2hw.tag_53.re;
  assign rcache_line[0][53].status_reg.status = reg2hw.status_53.q;//status_reg_t'(reg2hw.status_53.q);
  assign rcache_line[0][53].status_reg.qe    = reg2hw.status_53.qe;
  assign rcache_line[0][53].status_reg.re    = reg2hw.status_53.re;


  assign rcache_line[0][54].tag_reg.tag      = reg2hw.tag_54.q;
  assign rcache_line[0][54].tag_reg.qe       = reg2hw.tag_54.qe;
  assign rcache_line[0][54].tag_reg.re       = reg2hw.tag_54.re;
  assign rcache_line[0][54].status_reg.status = reg2hw.status_54.q;//status_reg_t'(reg2hw.status_54.q);
  assign rcache_line[0][54].status_reg.qe    = reg2hw.status_54.qe;
  assign rcache_line[0][54].status_reg.re    = reg2hw.status_54.re;


  assign rcache_line[0][55].tag_reg.tag      = reg2hw.tag_55.q;
  assign rcache_line[0][55].tag_reg.qe       = reg2hw.tag_55.qe;
  assign rcache_line[0][55].tag_reg.re       = reg2hw.tag_55.re;
  assign rcache_line[0][55].status_reg.status = reg2hw.status_55.q;//status_reg_t'(reg2hw.status_55.q);
  assign rcache_line[0][55].status_reg.qe    = reg2hw.status_55.qe;
  assign rcache_line[0][55].status_reg.re    = reg2hw.status_55.re;


  assign rcache_line[0][56].tag_reg.tag      = reg2hw.tag_56.q;
  assign rcache_line[0][56].tag_reg.qe       = reg2hw.tag_56.qe;
  assign rcache_line[0][56].tag_reg.re       = reg2hw.tag_56.re;
  assign rcache_line[0][56].status_reg.status = reg2hw.status_56.q;//status_reg_t'(reg2hw.status_56.q);
  assign rcache_line[0][56].status_reg.qe    = reg2hw.status_56.qe;
  assign rcache_line[0][56].status_reg.re    = reg2hw.status_56.re;


  assign rcache_line[0][57].tag_reg.tag      = reg2hw.tag_57.q;
  assign rcache_line[0][57].tag_reg.qe       = reg2hw.tag_57.qe;
  assign rcache_line[0][57].tag_reg.re       = reg2hw.tag_57.re;
  assign rcache_line[0][57].status_reg.status = reg2hw.status_57.q;//status_reg_t'(reg2hw.status_57.q);
  assign rcache_line[0][57].status_reg.qe    = reg2hw.status_57.qe;
  assign rcache_line[0][57].status_reg.re    = reg2hw.status_57.re;


  assign rcache_line[0][58].tag_reg.tag      = reg2hw.tag_58.q;
  assign rcache_line[0][58].tag_reg.qe       = reg2hw.tag_58.qe;
  assign rcache_line[0][58].tag_reg.re       = reg2hw.tag_58.re;
  assign rcache_line[0][58].status_reg.status = reg2hw.status_58.q;//status_reg_t'(reg2hw.status_58.q);
  assign rcache_line[0][58].status_reg.qe    = reg2hw.status_58.qe;
  assign rcache_line[0][58].status_reg.re    = reg2hw.status_58.re;


  assign rcache_line[0][59].tag_reg.tag      = reg2hw.tag_59.q;
  assign rcache_line[0][59].tag_reg.qe       = reg2hw.tag_59.qe;
  assign rcache_line[0][59].tag_reg.re       = reg2hw.tag_59.re;
  assign rcache_line[0][59].status_reg.status = reg2hw.status_59.q;//status_reg_t'(reg2hw.status_59.q);
  assign rcache_line[0][59].status_reg.qe    = reg2hw.status_59.qe;
  assign rcache_line[0][59].status_reg.re    = reg2hw.status_59.re;


  assign rcache_line[0][60].tag_reg.tag      = reg2hw.tag_60.q;
  assign rcache_line[0][60].tag_reg.qe       = reg2hw.tag_60.qe;
  assign rcache_line[0][60].tag_reg.re       = reg2hw.tag_60.re;
  assign rcache_line[0][60].status_reg.status = reg2hw.status_60.q;//status_reg_t'(reg2hw.status_60.q);
  assign rcache_line[0][60].status_reg.qe    = reg2hw.status_60.qe;
  assign rcache_line[0][60].status_reg.re    = reg2hw.status_60.re;


  assign rcache_line[0][61].tag_reg.tag      = reg2hw.tag_61.q;
  assign rcache_line[0][61].tag_reg.qe       = reg2hw.tag_61.qe;
  assign rcache_line[0][61].tag_reg.re       = reg2hw.tag_61.re;
  assign rcache_line[0][61].status_reg.status = reg2hw.status_61.q;//status_reg_t'(reg2hw.status_61.q);
  assign rcache_line[0][61].status_reg.qe    = reg2hw.status_61.qe;
  assign rcache_line[0][61].status_reg.re    = reg2hw.status_61.re;


  assign rcache_line[0][62].tag_reg.tag      = reg2hw.tag_62.q;
  assign rcache_line[0][62].tag_reg.qe       = reg2hw.tag_62.qe;
  assign rcache_line[0][62].tag_reg.re       = reg2hw.tag_62.re;
  assign rcache_line[0][62].status_reg.status = reg2hw.status_62.q;//status_reg_t'(reg2hw.status_62.q);
  assign rcache_line[0][62].status_reg.qe    = reg2hw.status_62.qe;
  assign rcache_line[0][62].status_reg.re    = reg2hw.status_62.re;


  assign rcache_line[0][63].tag_reg.tag      = reg2hw.tag_63.q;
  assign rcache_line[0][63].tag_reg.qe       = reg2hw.tag_63.qe;
  assign rcache_line[0][63].tag_reg.re       = reg2hw.tag_63.re;
  assign rcache_line[0][63].status_reg.status = reg2hw.status_63.q;//status_reg_t'(reg2hw.status_63.q);
  assign rcache_line[0][63].status_reg.qe    = reg2hw.status_63.qe;
  assign rcache_line[0][63].status_reg.re    = reg2hw.status_63.re;


  assign rcache_line[0][64].tag_reg.tag      = reg2hw.tag_64.q;
  assign rcache_line[0][64].tag_reg.qe       = reg2hw.tag_64.qe;
  assign rcache_line[0][64].tag_reg.re       = reg2hw.tag_64.re;
  assign rcache_line[0][64].status_reg.status = reg2hw.status_64.q;//status_reg_t'(reg2hw.status_64.q);
  assign rcache_line[0][64].status_reg.qe    = reg2hw.status_64.qe;
  assign rcache_line[0][64].status_reg.re    = reg2hw.status_64.re;


  assign rcache_line[0][65].tag_reg.tag      = reg2hw.tag_65.q;
  assign rcache_line[0][65].tag_reg.qe       = reg2hw.tag_65.qe;
  assign rcache_line[0][65].tag_reg.re       = reg2hw.tag_65.re;
  assign rcache_line[0][65].status_reg.status = reg2hw.status_65.q;//status_reg_t'(reg2hw.status_65.q);
  assign rcache_line[0][65].status_reg.qe    = reg2hw.status_65.qe;
  assign rcache_line[0][65].status_reg.re    = reg2hw.status_65.re;


  assign rcache_line[0][66].tag_reg.tag      = reg2hw.tag_66.q;
  assign rcache_line[0][66].tag_reg.qe       = reg2hw.tag_66.qe;
  assign rcache_line[0][66].tag_reg.re       = reg2hw.tag_66.re;
  assign rcache_line[0][66].status_reg.status = reg2hw.status_66.q;//status_reg_t'(reg2hw.status_66.q);
  assign rcache_line[0][66].status_reg.qe    = reg2hw.status_66.qe;
  assign rcache_line[0][66].status_reg.re    = reg2hw.status_66.re;


  assign rcache_line[0][67].tag_reg.tag      = reg2hw.tag_67.q;
  assign rcache_line[0][67].tag_reg.qe       = reg2hw.tag_67.qe;
  assign rcache_line[0][67].tag_reg.re       = reg2hw.tag_67.re;
  assign rcache_line[0][67].status_reg.status = reg2hw.status_67.q;//status_reg_t'(reg2hw.status_67.q);
  assign rcache_line[0][67].status_reg.qe    = reg2hw.status_67.qe;
  assign rcache_line[0][67].status_reg.re    = reg2hw.status_67.re;


  assign rcache_line[0][68].tag_reg.tag      = reg2hw.tag_68.q;
  assign rcache_line[0][68].tag_reg.qe       = reg2hw.tag_68.qe;
  assign rcache_line[0][68].tag_reg.re       = reg2hw.tag_68.re;
  assign rcache_line[0][68].status_reg.status = reg2hw.status_68.q;//status_reg_t'(reg2hw.status_68.q);
  assign rcache_line[0][68].status_reg.qe    = reg2hw.status_68.qe;
  assign rcache_line[0][68].status_reg.re    = reg2hw.status_68.re;


  assign rcache_line[0][69].tag_reg.tag      = reg2hw.tag_69.q;
  assign rcache_line[0][69].tag_reg.qe       = reg2hw.tag_69.qe;
  assign rcache_line[0][69].tag_reg.re       = reg2hw.tag_69.re;
  assign rcache_line[0][69].status_reg.status = reg2hw.status_69.q;//status_reg_t'(reg2hw.status_69.q);
  assign rcache_line[0][69].status_reg.qe    = reg2hw.status_69.qe;
  assign rcache_line[0][69].status_reg.re    = reg2hw.status_69.re;


  assign rcache_line[0][70].tag_reg.tag      = reg2hw.tag_70.q;
  assign rcache_line[0][70].tag_reg.qe       = reg2hw.tag_70.qe;
  assign rcache_line[0][70].tag_reg.re       = reg2hw.tag_70.re;
  assign rcache_line[0][70].status_reg.status = reg2hw.status_70.q;//status_reg_t'(reg2hw.status_70.q);
  assign rcache_line[0][70].status_reg.qe    = reg2hw.status_70.qe;
  assign rcache_line[0][70].status_reg.re    = reg2hw.status_70.re;


  assign rcache_line[0][71].tag_reg.tag      = reg2hw.tag_71.q;
  assign rcache_line[0][71].tag_reg.qe       = reg2hw.tag_71.qe;
  assign rcache_line[0][71].tag_reg.re       = reg2hw.tag_71.re;
  assign rcache_line[0][71].status_reg.status = reg2hw.status_71.q;//status_reg_t'(reg2hw.status_71.q);
  assign rcache_line[0][71].status_reg.qe    = reg2hw.status_71.qe;
  assign rcache_line[0][71].status_reg.re    = reg2hw.status_71.re;


  assign rcache_line[0][72].tag_reg.tag      = reg2hw.tag_72.q;
  assign rcache_line[0][72].tag_reg.qe       = reg2hw.tag_72.qe;
  assign rcache_line[0][72].tag_reg.re       = reg2hw.tag_72.re;
  assign rcache_line[0][72].status_reg.status = reg2hw.status_72.q;//status_reg_t'(reg2hw.status_72.q);
  assign rcache_line[0][72].status_reg.qe    = reg2hw.status_72.qe;
  assign rcache_line[0][72].status_reg.re    = reg2hw.status_72.re;


  assign rcache_line[0][73].tag_reg.tag      = reg2hw.tag_73.q;
  assign rcache_line[0][73].tag_reg.qe       = reg2hw.tag_73.qe;
  assign rcache_line[0][73].tag_reg.re       = reg2hw.tag_73.re;
  assign rcache_line[0][73].status_reg.status = reg2hw.status_73.q;//status_reg_t'(reg2hw.status_73.q);
  assign rcache_line[0][73].status_reg.qe    = reg2hw.status_73.qe;
  assign rcache_line[0][73].status_reg.re    = reg2hw.status_73.re;


  assign rcache_line[0][74].tag_reg.tag      = reg2hw.tag_74.q;
  assign rcache_line[0][74].tag_reg.qe       = reg2hw.tag_74.qe;
  assign rcache_line[0][74].tag_reg.re       = reg2hw.tag_74.re;
  assign rcache_line[0][74].status_reg.status = reg2hw.status_74.q;//status_reg_t'(reg2hw.status_74.q);
  assign rcache_line[0][74].status_reg.qe    = reg2hw.status_74.qe;
  assign rcache_line[0][74].status_reg.re    = reg2hw.status_74.re;


  assign rcache_line[0][75].tag_reg.tag      = reg2hw.tag_75.q;
  assign rcache_line[0][75].tag_reg.qe       = reg2hw.tag_75.qe;
  assign rcache_line[0][75].tag_reg.re       = reg2hw.tag_75.re;
  assign rcache_line[0][75].status_reg.status = reg2hw.status_75.q;//status_reg_t'(reg2hw.status_75.q);
  assign rcache_line[0][75].status_reg.qe    = reg2hw.status_75.qe;
  assign rcache_line[0][75].status_reg.re    = reg2hw.status_75.re;


  assign rcache_line[0][76].tag_reg.tag      = reg2hw.tag_76.q;
  assign rcache_line[0][76].tag_reg.qe       = reg2hw.tag_76.qe;
  assign rcache_line[0][76].tag_reg.re       = reg2hw.tag_76.re;
  assign rcache_line[0][76].status_reg.status = reg2hw.status_76.q;//status_reg_t'(reg2hw.status_76.q);
  assign rcache_line[0][76].status_reg.qe    = reg2hw.status_76.qe;
  assign rcache_line[0][76].status_reg.re    = reg2hw.status_76.re;


  assign rcache_line[0][77].tag_reg.tag      = reg2hw.tag_77.q;
  assign rcache_line[0][77].tag_reg.qe       = reg2hw.tag_77.qe;
  assign rcache_line[0][77].tag_reg.re       = reg2hw.tag_77.re;
  assign rcache_line[0][77].status_reg.status = reg2hw.status_77.q;//status_reg_t'(reg2hw.status_77.q);
  assign rcache_line[0][77].status_reg.qe    = reg2hw.status_77.qe;
  assign rcache_line[0][77].status_reg.re    = reg2hw.status_77.re;


  assign rcache_line[0][78].tag_reg.tag      = reg2hw.tag_78.q;
  assign rcache_line[0][78].tag_reg.qe       = reg2hw.tag_78.qe;
  assign rcache_line[0][78].tag_reg.re       = reg2hw.tag_78.re;
  assign rcache_line[0][78].status_reg.status = reg2hw.status_78.q;//status_reg_t'(reg2hw.status_78.q);
  assign rcache_line[0][78].status_reg.qe    = reg2hw.status_78.qe;
  assign rcache_line[0][78].status_reg.re    = reg2hw.status_78.re;


  assign rcache_line[0][79].tag_reg.tag      = reg2hw.tag_79.q;
  assign rcache_line[0][79].tag_reg.qe       = reg2hw.tag_79.qe;
  assign rcache_line[0][79].tag_reg.re       = reg2hw.tag_79.re;
  assign rcache_line[0][79].status_reg.status = reg2hw.status_79.q;//status_reg_t'(reg2hw.status_79.q);
  assign rcache_line[0][79].status_reg.qe    = reg2hw.status_79.qe;
  assign rcache_line[0][79].status_reg.re    = reg2hw.status_79.re;


  assign rcache_line[0][80].tag_reg.tag      = reg2hw.tag_80.q;
  assign rcache_line[0][80].tag_reg.qe       = reg2hw.tag_80.qe;
  assign rcache_line[0][80].tag_reg.re       = reg2hw.tag_80.re;
  assign rcache_line[0][80].status_reg.status = reg2hw.status_80.q;//status_reg_t'(reg2hw.status_80.q);
  assign rcache_line[0][80].status_reg.qe    = reg2hw.status_80.qe;
  assign rcache_line[0][80].status_reg.re    = reg2hw.status_80.re;


  assign rcache_line[0][81].tag_reg.tag      = reg2hw.tag_81.q;
  assign rcache_line[0][81].tag_reg.qe       = reg2hw.tag_81.qe;
  assign rcache_line[0][81].tag_reg.re       = reg2hw.tag_81.re;
  assign rcache_line[0][81].status_reg.status = reg2hw.status_81.q;//status_reg_t'(reg2hw.status_81.q);
  assign rcache_line[0][81].status_reg.qe    = reg2hw.status_81.qe;
  assign rcache_line[0][81].status_reg.re    = reg2hw.status_81.re;


  assign rcache_line[0][82].tag_reg.tag      = reg2hw.tag_82.q;
  assign rcache_line[0][82].tag_reg.qe       = reg2hw.tag_82.qe;
  assign rcache_line[0][82].tag_reg.re       = reg2hw.tag_82.re;
  assign rcache_line[0][82].status_reg.status = reg2hw.status_82.q;//status_reg_t'(reg2hw.status_82.q);
  assign rcache_line[0][82].status_reg.qe    = reg2hw.status_82.qe;
  assign rcache_line[0][82].status_reg.re    = reg2hw.status_82.re;


  assign rcache_line[0][83].tag_reg.tag      = reg2hw.tag_83.q;
  assign rcache_line[0][83].tag_reg.qe       = reg2hw.tag_83.qe;
  assign rcache_line[0][83].tag_reg.re       = reg2hw.tag_83.re;
  assign rcache_line[0][83].status_reg.status = reg2hw.status_83.q;//status_reg_t'(reg2hw.status_83.q);
  assign rcache_line[0][83].status_reg.qe    = reg2hw.status_83.qe;
  assign rcache_line[0][83].status_reg.re    = reg2hw.status_83.re;


  assign rcache_line[0][84].tag_reg.tag      = reg2hw.tag_84.q;
  assign rcache_line[0][84].tag_reg.qe       = reg2hw.tag_84.qe;
  assign rcache_line[0][84].tag_reg.re       = reg2hw.tag_84.re;
  assign rcache_line[0][84].status_reg.status = reg2hw.status_84.q;//status_reg_t'(reg2hw.status_84.q);
  assign rcache_line[0][84].status_reg.qe    = reg2hw.status_84.qe;
  assign rcache_line[0][84].status_reg.re    = reg2hw.status_84.re;


  assign rcache_line[0][85].tag_reg.tag      = reg2hw.tag_85.q;
  assign rcache_line[0][85].tag_reg.qe       = reg2hw.tag_85.qe;
  assign rcache_line[0][85].tag_reg.re       = reg2hw.tag_85.re;
  assign rcache_line[0][85].status_reg.status = reg2hw.status_85.q;//status_reg_t'(reg2hw.status_85.q);
  assign rcache_line[0][85].status_reg.qe    = reg2hw.status_85.qe;
  assign rcache_line[0][85].status_reg.re    = reg2hw.status_85.re;


  assign rcache_line[0][86].tag_reg.tag      = reg2hw.tag_86.q;
  assign rcache_line[0][86].tag_reg.qe       = reg2hw.tag_86.qe;
  assign rcache_line[0][86].tag_reg.re       = reg2hw.tag_86.re;
  assign rcache_line[0][86].status_reg.status = reg2hw.status_86.q;//status_reg_t'(reg2hw.status_86.q);
  assign rcache_line[0][86].status_reg.qe    = reg2hw.status_86.qe;
  assign rcache_line[0][86].status_reg.re    = reg2hw.status_86.re;


  assign rcache_line[0][87].tag_reg.tag      = reg2hw.tag_87.q;
  assign rcache_line[0][87].tag_reg.qe       = reg2hw.tag_87.qe;
  assign rcache_line[0][87].tag_reg.re       = reg2hw.tag_87.re;
  assign rcache_line[0][87].status_reg.status = reg2hw.status_87.q;//status_reg_t'(reg2hw.status_87.q);
  assign rcache_line[0][87].status_reg.qe    = reg2hw.status_87.qe;
  assign rcache_line[0][87].status_reg.re    = reg2hw.status_87.re;


  assign rcache_line[0][88].tag_reg.tag      = reg2hw.tag_88.q;
  assign rcache_line[0][88].tag_reg.qe       = reg2hw.tag_88.qe;
  assign rcache_line[0][88].tag_reg.re       = reg2hw.tag_88.re;
  assign rcache_line[0][88].status_reg.status = reg2hw.status_88.q;//status_reg_t'(reg2hw.status_88.q);
  assign rcache_line[0][88].status_reg.qe    = reg2hw.status_88.qe;
  assign rcache_line[0][88].status_reg.re    = reg2hw.status_88.re;


  assign rcache_line[0][89].tag_reg.tag      = reg2hw.tag_89.q;
  assign rcache_line[0][89].tag_reg.qe       = reg2hw.tag_89.qe;
  assign rcache_line[0][89].tag_reg.re       = reg2hw.tag_89.re;
  assign rcache_line[0][89].status_reg.status = reg2hw.status_89.q;//status_reg_t'(reg2hw.status_89.q);
  assign rcache_line[0][89].status_reg.qe    = reg2hw.status_89.qe;
  assign rcache_line[0][89].status_reg.re    = reg2hw.status_89.re;


  assign rcache_line[0][90].tag_reg.tag      = reg2hw.tag_90.q;
  assign rcache_line[0][90].tag_reg.qe       = reg2hw.tag_90.qe;
  assign rcache_line[0][90].tag_reg.re       = reg2hw.tag_90.re;
  assign rcache_line[0][90].status_reg.status = reg2hw.status_90.q;//status_reg_t'(reg2hw.status_90.q);
  assign rcache_line[0][90].status_reg.qe    = reg2hw.status_90.qe;
  assign rcache_line[0][90].status_reg.re    = reg2hw.status_90.re;


  assign rcache_line[0][91].tag_reg.tag      = reg2hw.tag_91.q;
  assign rcache_line[0][91].tag_reg.qe       = reg2hw.tag_91.qe;
  assign rcache_line[0][91].tag_reg.re       = reg2hw.tag_91.re;
  assign rcache_line[0][91].status_reg.status = reg2hw.status_91.q;//status_reg_t'(reg2hw.status_91.q);
  assign rcache_line[0][91].status_reg.qe    = reg2hw.status_91.qe;
  assign rcache_line[0][91].status_reg.re    = reg2hw.status_91.re;


  assign rcache_line[0][92].tag_reg.tag      = reg2hw.tag_92.q;
  assign rcache_line[0][92].tag_reg.qe       = reg2hw.tag_92.qe;
  assign rcache_line[0][92].tag_reg.re       = reg2hw.tag_92.re;
  assign rcache_line[0][92].status_reg.status = reg2hw.status_92.q;//status_reg_t'(reg2hw.status_92.q);
  assign rcache_line[0][92].status_reg.qe    = reg2hw.status_92.qe;
  assign rcache_line[0][92].status_reg.re    = reg2hw.status_92.re;


  assign rcache_line[0][93].tag_reg.tag      = reg2hw.tag_93.q;
  assign rcache_line[0][93].tag_reg.qe       = reg2hw.tag_93.qe;
  assign rcache_line[0][93].tag_reg.re       = reg2hw.tag_93.re;
  assign rcache_line[0][93].status_reg.status = reg2hw.status_93.q;//status_reg_t'(reg2hw.status_93.q);
  assign rcache_line[0][93].status_reg.qe    = reg2hw.status_93.qe;
  assign rcache_line[0][93].status_reg.re    = reg2hw.status_93.re;


  assign rcache_line[0][94].tag_reg.tag      = reg2hw.tag_94.q;
  assign rcache_line[0][94].tag_reg.qe       = reg2hw.tag_94.qe;
  assign rcache_line[0][94].tag_reg.re       = reg2hw.tag_94.re;
  assign rcache_line[0][94].status_reg.status = reg2hw.status_94.q;//status_reg_t'(reg2hw.status_94.q);
  assign rcache_line[0][94].status_reg.qe    = reg2hw.status_94.qe;
  assign rcache_line[0][94].status_reg.re    = reg2hw.status_94.re;


  assign rcache_line[0][95].tag_reg.tag      = reg2hw.tag_95.q;
  assign rcache_line[0][95].tag_reg.qe       = reg2hw.tag_95.qe;
  assign rcache_line[0][95].tag_reg.re       = reg2hw.tag_95.re;
  assign rcache_line[0][95].status_reg.status = reg2hw.status_95.q;//status_reg_t'(reg2hw.status_95.q);
  assign rcache_line[0][95].status_reg.qe    = reg2hw.status_95.qe;
  assign rcache_line[0][95].status_reg.re    = reg2hw.status_95.re;


  assign rcache_line[0][96].tag_reg.tag      = reg2hw.tag_96.q;
  assign rcache_line[0][96].tag_reg.qe       = reg2hw.tag_96.qe;
  assign rcache_line[0][96].tag_reg.re       = reg2hw.tag_96.re;
  assign rcache_line[0][96].status_reg.status = reg2hw.status_96.q;//status_reg_t'(reg2hw.status_96.q);
  assign rcache_line[0][96].status_reg.qe    = reg2hw.status_96.qe;
  assign rcache_line[0][96].status_reg.re    = reg2hw.status_96.re;


  assign rcache_line[0][97].tag_reg.tag      = reg2hw.tag_97.q;
  assign rcache_line[0][97].tag_reg.qe       = reg2hw.tag_97.qe;
  assign rcache_line[0][97].tag_reg.re       = reg2hw.tag_97.re;
  assign rcache_line[0][97].status_reg.status = reg2hw.status_97.q;//status_reg_t'(reg2hw.status_97.q);
  assign rcache_line[0][97].status_reg.qe    = reg2hw.status_97.qe;
  assign rcache_line[0][97].status_reg.re    = reg2hw.status_97.re;


  assign rcache_line[0][98].tag_reg.tag      = reg2hw.tag_98.q;
  assign rcache_line[0][98].tag_reg.qe       = reg2hw.tag_98.qe;
  assign rcache_line[0][98].tag_reg.re       = reg2hw.tag_98.re;
  assign rcache_line[0][98].status_reg.status = reg2hw.status_98.q;//status_reg_t'(reg2hw.status_98.q);
  assign rcache_line[0][98].status_reg.qe    = reg2hw.status_98.qe;
  assign rcache_line[0][98].status_reg.re    = reg2hw.status_98.re;


  assign rcache_line[0][99].tag_reg.tag      = reg2hw.tag_99.q;
  assign rcache_line[0][99].tag_reg.qe       = reg2hw.tag_99.qe;
  assign rcache_line[0][99].tag_reg.re       = reg2hw.tag_99.re;
  assign rcache_line[0][99].status_reg.status = reg2hw.status_99.q;//status_reg_t'(reg2hw.status_99.q);
  assign rcache_line[0][99].status_reg.qe    = reg2hw.status_99.qe;
  assign rcache_line[0][99].status_reg.re    = reg2hw.status_99.re;


  assign rcache_line[0][100].tag_reg.tag      = reg2hw.tag_100.q;
  assign rcache_line[0][100].tag_reg.qe       = reg2hw.tag_100.qe;
  assign rcache_line[0][100].tag_reg.re       = reg2hw.tag_100.re;
  assign rcache_line[0][100].status_reg.status = reg2hw.status_100.q;//status_reg_t'(reg2hw.status_100.q);
  assign rcache_line[0][100].status_reg.qe    = reg2hw.status_100.qe;
  assign rcache_line[0][100].status_reg.re    = reg2hw.status_100.re;


  assign rcache_line[0][101].tag_reg.tag      = reg2hw.tag_101.q;
  assign rcache_line[0][101].tag_reg.qe       = reg2hw.tag_101.qe;
  assign rcache_line[0][101].tag_reg.re       = reg2hw.tag_101.re;
  assign rcache_line[0][101].status_reg.status = reg2hw.status_101.q;//status_reg_t'(reg2hw.status_101.q);
  assign rcache_line[0][101].status_reg.qe    = reg2hw.status_101.qe;
  assign rcache_line[0][101].status_reg.re    = reg2hw.status_101.re;


  assign rcache_line[0][102].tag_reg.tag      = reg2hw.tag_102.q;
  assign rcache_line[0][102].tag_reg.qe       = reg2hw.tag_102.qe;
  assign rcache_line[0][102].tag_reg.re       = reg2hw.tag_102.re;
  assign rcache_line[0][102].status_reg.status = reg2hw.status_102.q;//status_reg_t'(reg2hw.status_102.q);
  assign rcache_line[0][102].status_reg.qe    = reg2hw.status_102.qe;
  assign rcache_line[0][102].status_reg.re    = reg2hw.status_102.re;


  assign rcache_line[0][103].tag_reg.tag      = reg2hw.tag_103.q;
  assign rcache_line[0][103].tag_reg.qe       = reg2hw.tag_103.qe;
  assign rcache_line[0][103].tag_reg.re       = reg2hw.tag_103.re;
  assign rcache_line[0][103].status_reg.status = reg2hw.status_103.q;//status_reg_t'(reg2hw.status_103.q);
  assign rcache_line[0][103].status_reg.qe    = reg2hw.status_103.qe;
  assign rcache_line[0][103].status_reg.re    = reg2hw.status_103.re;


  assign rcache_line[0][104].tag_reg.tag      = reg2hw.tag_104.q;
  assign rcache_line[0][104].tag_reg.qe       = reg2hw.tag_104.qe;
  assign rcache_line[0][104].tag_reg.re       = reg2hw.tag_104.re;
  assign rcache_line[0][104].status_reg.status = reg2hw.status_104.q;//status_reg_t'(reg2hw.status_104.q);
  assign rcache_line[0][104].status_reg.qe    = reg2hw.status_104.qe;
  assign rcache_line[0][104].status_reg.re    = reg2hw.status_104.re;


  assign rcache_line[0][105].tag_reg.tag      = reg2hw.tag_105.q;
  assign rcache_line[0][105].tag_reg.qe       = reg2hw.tag_105.qe;
  assign rcache_line[0][105].tag_reg.re       = reg2hw.tag_105.re;
  assign rcache_line[0][105].status_reg.status = reg2hw.status_105.q;//status_reg_t'(reg2hw.status_105.q);
  assign rcache_line[0][105].status_reg.qe    = reg2hw.status_105.qe;
  assign rcache_line[0][105].status_reg.re    = reg2hw.status_105.re;


  assign rcache_line[0][106].tag_reg.tag      = reg2hw.tag_106.q;
  assign rcache_line[0][106].tag_reg.qe       = reg2hw.tag_106.qe;
  assign rcache_line[0][106].tag_reg.re       = reg2hw.tag_106.re;
  assign rcache_line[0][106].status_reg.status = reg2hw.status_106.q;//status_reg_t'(reg2hw.status_106.q);
  assign rcache_line[0][106].status_reg.qe    = reg2hw.status_106.qe;
  assign rcache_line[0][106].status_reg.re    = reg2hw.status_106.re;


  assign rcache_line[0][107].tag_reg.tag      = reg2hw.tag_107.q;
  assign rcache_line[0][107].tag_reg.qe       = reg2hw.tag_107.qe;
  assign rcache_line[0][107].tag_reg.re       = reg2hw.tag_107.re;
  assign rcache_line[0][107].status_reg.status = reg2hw.status_107.q;//status_reg_t'(reg2hw.status_107.q);
  assign rcache_line[0][107].status_reg.qe    = reg2hw.status_107.qe;
  assign rcache_line[0][107].status_reg.re    = reg2hw.status_107.re;


  assign rcache_line[0][108].tag_reg.tag      = reg2hw.tag_108.q;
  assign rcache_line[0][108].tag_reg.qe       = reg2hw.tag_108.qe;
  assign rcache_line[0][108].tag_reg.re       = reg2hw.tag_108.re;
  assign rcache_line[0][108].status_reg.status = reg2hw.status_108.q;//status_reg_t'(reg2hw.status_108.q);
  assign rcache_line[0][108].status_reg.qe    = reg2hw.status_108.qe;
  assign rcache_line[0][108].status_reg.re    = reg2hw.status_108.re;


  assign rcache_line[0][109].tag_reg.tag      = reg2hw.tag_109.q;
  assign rcache_line[0][109].tag_reg.qe       = reg2hw.tag_109.qe;
  assign rcache_line[0][109].tag_reg.re       = reg2hw.tag_109.re;
  assign rcache_line[0][109].status_reg.status = reg2hw.status_109.q;//status_reg_t'(reg2hw.status_109.q);
  assign rcache_line[0][109].status_reg.qe    = reg2hw.status_109.qe;
  assign rcache_line[0][109].status_reg.re    = reg2hw.status_109.re;


  assign rcache_line[0][110].tag_reg.tag      = reg2hw.tag_110.q;
  assign rcache_line[0][110].tag_reg.qe       = reg2hw.tag_110.qe;
  assign rcache_line[0][110].tag_reg.re       = reg2hw.tag_110.re;
  assign rcache_line[0][110].status_reg.status = reg2hw.status_110.q;//status_reg_t'(reg2hw.status_110.q);
  assign rcache_line[0][110].status_reg.qe    = reg2hw.status_110.qe;
  assign rcache_line[0][110].status_reg.re    = reg2hw.status_110.re;


  assign rcache_line[0][111].tag_reg.tag      = reg2hw.tag_111.q;
  assign rcache_line[0][111].tag_reg.qe       = reg2hw.tag_111.qe;
  assign rcache_line[0][111].tag_reg.re       = reg2hw.tag_111.re;
  assign rcache_line[0][111].status_reg.status = reg2hw.status_111.q;//status_reg_t'(reg2hw.status_111.q);
  assign rcache_line[0][111].status_reg.qe    = reg2hw.status_111.qe;
  assign rcache_line[0][111].status_reg.re    = reg2hw.status_111.re;


  assign rcache_line[0][112].tag_reg.tag      = reg2hw.tag_112.q;
  assign rcache_line[0][112].tag_reg.qe       = reg2hw.tag_112.qe;
  assign rcache_line[0][112].tag_reg.re       = reg2hw.tag_112.re;
  assign rcache_line[0][112].status_reg.status = reg2hw.status_112.q;//status_reg_t'(reg2hw.status_112.q);
  assign rcache_line[0][112].status_reg.qe    = reg2hw.status_112.qe;
  assign rcache_line[0][112].status_reg.re    = reg2hw.status_112.re;


  assign rcache_line[0][113].tag_reg.tag      = reg2hw.tag_113.q;
  assign rcache_line[0][113].tag_reg.qe       = reg2hw.tag_113.qe;
  assign rcache_line[0][113].tag_reg.re       = reg2hw.tag_113.re;
  assign rcache_line[0][113].status_reg.status = reg2hw.status_113.q;//status_reg_t'(reg2hw.status_113.q);
  assign rcache_line[0][113].status_reg.qe    = reg2hw.status_113.qe;
  assign rcache_line[0][113].status_reg.re    = reg2hw.status_113.re;


  assign rcache_line[0][114].tag_reg.tag      = reg2hw.tag_114.q;
  assign rcache_line[0][114].tag_reg.qe       = reg2hw.tag_114.qe;
  assign rcache_line[0][114].tag_reg.re       = reg2hw.tag_114.re;
  assign rcache_line[0][114].status_reg.status = reg2hw.status_114.q;//status_reg_t'(reg2hw.status_114.q);
  assign rcache_line[0][114].status_reg.qe    = reg2hw.status_114.qe;
  assign rcache_line[0][114].status_reg.re    = reg2hw.status_114.re;


  assign rcache_line[0][115].tag_reg.tag      = reg2hw.tag_115.q;
  assign rcache_line[0][115].tag_reg.qe       = reg2hw.tag_115.qe;
  assign rcache_line[0][115].tag_reg.re       = reg2hw.tag_115.re;
  assign rcache_line[0][115].status_reg.status = reg2hw.status_115.q;//status_reg_t'(reg2hw.status_115.q);
  assign rcache_line[0][115].status_reg.qe    = reg2hw.status_115.qe;
  assign rcache_line[0][115].status_reg.re    = reg2hw.status_115.re;


  assign rcache_line[0][116].tag_reg.tag      = reg2hw.tag_116.q;
  assign rcache_line[0][116].tag_reg.qe       = reg2hw.tag_116.qe;
  assign rcache_line[0][116].tag_reg.re       = reg2hw.tag_116.re;
  assign rcache_line[0][116].status_reg.status = reg2hw.status_116.q;//status_reg_t'(reg2hw.status_116.q);
  assign rcache_line[0][116].status_reg.qe    = reg2hw.status_116.qe;
  assign rcache_line[0][116].status_reg.re    = reg2hw.status_116.re;


  assign rcache_line[0][117].tag_reg.tag      = reg2hw.tag_117.q;
  assign rcache_line[0][117].tag_reg.qe       = reg2hw.tag_117.qe;
  assign rcache_line[0][117].tag_reg.re       = reg2hw.tag_117.re;
  assign rcache_line[0][117].status_reg.status = reg2hw.status_117.q;//status_reg_t'(reg2hw.status_117.q);
  assign rcache_line[0][117].status_reg.qe    = reg2hw.status_117.qe;
  assign rcache_line[0][117].status_reg.re    = reg2hw.status_117.re;


  assign rcache_line[0][118].tag_reg.tag      = reg2hw.tag_118.q;
  assign rcache_line[0][118].tag_reg.qe       = reg2hw.tag_118.qe;
  assign rcache_line[0][118].tag_reg.re       = reg2hw.tag_118.re;
  assign rcache_line[0][118].status_reg.status = reg2hw.status_118.q;//status_reg_t'(reg2hw.status_118.q);
  assign rcache_line[0][118].status_reg.qe    = reg2hw.status_118.qe;
  assign rcache_line[0][118].status_reg.re    = reg2hw.status_118.re;


  assign rcache_line[0][119].tag_reg.tag      = reg2hw.tag_119.q;
  assign rcache_line[0][119].tag_reg.qe       = reg2hw.tag_119.qe;
  assign rcache_line[0][119].tag_reg.re       = reg2hw.tag_119.re;
  assign rcache_line[0][119].status_reg.status = reg2hw.status_119.q;//status_reg_t'(reg2hw.status_119.q);
  assign rcache_line[0][119].status_reg.qe    = reg2hw.status_119.qe;
  assign rcache_line[0][119].status_reg.re    = reg2hw.status_119.re;


  assign rcache_line[0][120].tag_reg.tag      = reg2hw.tag_120.q;
  assign rcache_line[0][120].tag_reg.qe       = reg2hw.tag_120.qe;
  assign rcache_line[0][120].tag_reg.re       = reg2hw.tag_120.re;
  assign rcache_line[0][120].status_reg.status = reg2hw.status_120.q;//status_reg_t'(reg2hw.status_120.q);
  assign rcache_line[0][120].status_reg.qe    = reg2hw.status_120.qe;
  assign rcache_line[0][120].status_reg.re    = reg2hw.status_120.re;


  assign rcache_line[0][121].tag_reg.tag      = reg2hw.tag_121.q;
  assign rcache_line[0][121].tag_reg.qe       = reg2hw.tag_121.qe;
  assign rcache_line[0][121].tag_reg.re       = reg2hw.tag_121.re;
  assign rcache_line[0][121].status_reg.status = reg2hw.status_121.q;//status_reg_t'(reg2hw.status_121.q);
  assign rcache_line[0][121].status_reg.qe    = reg2hw.status_121.qe;
  assign rcache_line[0][121].status_reg.re    = reg2hw.status_121.re;


  assign rcache_line[0][122].tag_reg.tag      = reg2hw.tag_122.q;
  assign rcache_line[0][122].tag_reg.qe       = reg2hw.tag_122.qe;
  assign rcache_line[0][122].tag_reg.re       = reg2hw.tag_122.re;
  assign rcache_line[0][122].status_reg.status = reg2hw.status_122.q;//status_reg_t'(reg2hw.status_122.q);
  assign rcache_line[0][122].status_reg.qe    = reg2hw.status_122.qe;
  assign rcache_line[0][122].status_reg.re    = reg2hw.status_122.re;


  assign rcache_line[0][123].tag_reg.tag      = reg2hw.tag_123.q;
  assign rcache_line[0][123].tag_reg.qe       = reg2hw.tag_123.qe;
  assign rcache_line[0][123].tag_reg.re       = reg2hw.tag_123.re;
  assign rcache_line[0][123].status_reg.status = reg2hw.status_123.q;//status_reg_t'(reg2hw.status_123.q);
  assign rcache_line[0][123].status_reg.qe    = reg2hw.status_123.qe;
  assign rcache_line[0][123].status_reg.re    = reg2hw.status_123.re;


  assign rcache_line[0][124].tag_reg.tag      = reg2hw.tag_124.q;
  assign rcache_line[0][124].tag_reg.qe       = reg2hw.tag_124.qe;
  assign rcache_line[0][124].tag_reg.re       = reg2hw.tag_124.re;
  assign rcache_line[0][124].status_reg.status = reg2hw.status_124.q;//status_reg_t'(reg2hw.status_124.q);
  assign rcache_line[0][124].status_reg.qe    = reg2hw.status_124.qe;
  assign rcache_line[0][124].status_reg.re    = reg2hw.status_124.re;


  assign rcache_line[0][125].tag_reg.tag      = reg2hw.tag_125.q;
  assign rcache_line[0][125].tag_reg.qe       = reg2hw.tag_125.qe;
  assign rcache_line[0][125].tag_reg.re       = reg2hw.tag_125.re;
  assign rcache_line[0][125].status_reg.status = reg2hw.status_125.q;//status_reg_t'(reg2hw.status_125.q);
  assign rcache_line[0][125].status_reg.qe    = reg2hw.status_125.qe;
  assign rcache_line[0][125].status_reg.re    = reg2hw.status_125.re;


  assign rcache_line[0][126].tag_reg.tag      = reg2hw.tag_126.q;
  assign rcache_line[0][126].tag_reg.qe       = reg2hw.tag_126.qe;
  assign rcache_line[0][126].tag_reg.re       = reg2hw.tag_126.re;
  assign rcache_line[0][126].status_reg.status = reg2hw.status_126.q;//status_reg_t'(reg2hw.status_126.q);
  assign rcache_line[0][126].status_reg.qe    = reg2hw.status_126.qe;
  assign rcache_line[0][126].status_reg.re    = reg2hw.status_126.re;


  assign rcache_line[0][127].tag_reg.tag      = reg2hw.tag_127.q;
  assign rcache_line[0][127].tag_reg.qe       = reg2hw.tag_127.qe;
  assign rcache_line[0][127].tag_reg.re       = reg2hw.tag_127.re;
  assign rcache_line[0][127].status_reg.status = reg2hw.status_127.q;//status_reg_t'(reg2hw.status_127.q);
  assign rcache_line[0][127].status_reg.qe    = reg2hw.status_127.qe;
  assign rcache_line[0][127].status_reg.re    = reg2hw.status_127.re;


  assign rcache_line[0][128].tag_reg.tag      = reg2hw.tag_128.q;
  assign rcache_line[0][128].tag_reg.qe       = reg2hw.tag_128.qe;
  assign rcache_line[0][128].tag_reg.re       = reg2hw.tag_128.re;
  assign rcache_line[0][128].status_reg.status = reg2hw.status_128.q;//status_reg_t'(reg2hw.status_128.q);
  assign rcache_line[0][128].status_reg.qe    = reg2hw.status_128.qe;
  assign rcache_line[0][128].status_reg.re    = reg2hw.status_128.re;


  assign rcache_line[0][129].tag_reg.tag      = reg2hw.tag_129.q;
  assign rcache_line[0][129].tag_reg.qe       = reg2hw.tag_129.qe;
  assign rcache_line[0][129].tag_reg.re       = reg2hw.tag_129.re;
  assign rcache_line[0][129].status_reg.status = reg2hw.status_129.q;//status_reg_t'(reg2hw.status_129.q);
  assign rcache_line[0][129].status_reg.qe    = reg2hw.status_129.qe;
  assign rcache_line[0][129].status_reg.re    = reg2hw.status_129.re;


  assign rcache_line[0][130].tag_reg.tag      = reg2hw.tag_130.q;
  assign rcache_line[0][130].tag_reg.qe       = reg2hw.tag_130.qe;
  assign rcache_line[0][130].tag_reg.re       = reg2hw.tag_130.re;
  assign rcache_line[0][130].status_reg.status = reg2hw.status_130.q;//status_reg_t'(reg2hw.status_130.q);
  assign rcache_line[0][130].status_reg.qe    = reg2hw.status_130.qe;
  assign rcache_line[0][130].status_reg.re    = reg2hw.status_130.re;


  assign rcache_line[0][131].tag_reg.tag      = reg2hw.tag_131.q;
  assign rcache_line[0][131].tag_reg.qe       = reg2hw.tag_131.qe;
  assign rcache_line[0][131].tag_reg.re       = reg2hw.tag_131.re;
  assign rcache_line[0][131].status_reg.status = reg2hw.status_131.q;//status_reg_t'(reg2hw.status_131.q);
  assign rcache_line[0][131].status_reg.qe    = reg2hw.status_131.qe;
  assign rcache_line[0][131].status_reg.re    = reg2hw.status_131.re;


  assign rcache_line[0][132].tag_reg.tag      = reg2hw.tag_132.q;
  assign rcache_line[0][132].tag_reg.qe       = reg2hw.tag_132.qe;
  assign rcache_line[0][132].tag_reg.re       = reg2hw.tag_132.re;
  assign rcache_line[0][132].status_reg.status = reg2hw.status_132.q;//status_reg_t'(reg2hw.status_132.q);
  assign rcache_line[0][132].status_reg.qe    = reg2hw.status_132.qe;
  assign rcache_line[0][132].status_reg.re    = reg2hw.status_132.re;


  assign rcache_line[0][133].tag_reg.tag      = reg2hw.tag_133.q;
  assign rcache_line[0][133].tag_reg.qe       = reg2hw.tag_133.qe;
  assign rcache_line[0][133].tag_reg.re       = reg2hw.tag_133.re;
  assign rcache_line[0][133].status_reg.status = reg2hw.status_133.q;//status_reg_t'(reg2hw.status_133.q);
  assign rcache_line[0][133].status_reg.qe    = reg2hw.status_133.qe;
  assign rcache_line[0][133].status_reg.re    = reg2hw.status_133.re;


  assign rcache_line[0][134].tag_reg.tag      = reg2hw.tag_134.q;
  assign rcache_line[0][134].tag_reg.qe       = reg2hw.tag_134.qe;
  assign rcache_line[0][134].tag_reg.re       = reg2hw.tag_134.re;
  assign rcache_line[0][134].status_reg.status = reg2hw.status_134.q;//status_reg_t'(reg2hw.status_134.q);
  assign rcache_line[0][134].status_reg.qe    = reg2hw.status_134.qe;
  assign rcache_line[0][134].status_reg.re    = reg2hw.status_134.re;


  assign rcache_line[0][135].tag_reg.tag      = reg2hw.tag_135.q;
  assign rcache_line[0][135].tag_reg.qe       = reg2hw.tag_135.qe;
  assign rcache_line[0][135].tag_reg.re       = reg2hw.tag_135.re;
  assign rcache_line[0][135].status_reg.status = reg2hw.status_135.q;//status_reg_t'(reg2hw.status_135.q);
  assign rcache_line[0][135].status_reg.qe    = reg2hw.status_135.qe;
  assign rcache_line[0][135].status_reg.re    = reg2hw.status_135.re;


  assign rcache_line[0][136].tag_reg.tag      = reg2hw.tag_136.q;
  assign rcache_line[0][136].tag_reg.qe       = reg2hw.tag_136.qe;
  assign rcache_line[0][136].tag_reg.re       = reg2hw.tag_136.re;
  assign rcache_line[0][136].status_reg.status = reg2hw.status_136.q;//status_reg_t'(reg2hw.status_136.q);
  assign rcache_line[0][136].status_reg.qe    = reg2hw.status_136.qe;
  assign rcache_line[0][136].status_reg.re    = reg2hw.status_136.re;


  assign rcache_line[0][137].tag_reg.tag      = reg2hw.tag_137.q;
  assign rcache_line[0][137].tag_reg.qe       = reg2hw.tag_137.qe;
  assign rcache_line[0][137].tag_reg.re       = reg2hw.tag_137.re;
  assign rcache_line[0][137].status_reg.status = reg2hw.status_137.q;//status_reg_t'(reg2hw.status_137.q);
  assign rcache_line[0][137].status_reg.qe    = reg2hw.status_137.qe;
  assign rcache_line[0][137].status_reg.re    = reg2hw.status_137.re;


  assign rcache_line[0][138].tag_reg.tag      = reg2hw.tag_138.q;
  assign rcache_line[0][138].tag_reg.qe       = reg2hw.tag_138.qe;
  assign rcache_line[0][138].tag_reg.re       = reg2hw.tag_138.re;
  assign rcache_line[0][138].status_reg.status = reg2hw.status_138.q;//status_reg_t'(reg2hw.status_138.q);
  assign rcache_line[0][138].status_reg.qe    = reg2hw.status_138.qe;
  assign rcache_line[0][138].status_reg.re    = reg2hw.status_138.re;


  assign rcache_line[0][139].tag_reg.tag      = reg2hw.tag_139.q;
  assign rcache_line[0][139].tag_reg.qe       = reg2hw.tag_139.qe;
  assign rcache_line[0][139].tag_reg.re       = reg2hw.tag_139.re;
  assign rcache_line[0][139].status_reg.status = reg2hw.status_139.q;//status_reg_t'(reg2hw.status_139.q);
  assign rcache_line[0][139].status_reg.qe    = reg2hw.status_139.qe;
  assign rcache_line[0][139].status_reg.re    = reg2hw.status_139.re;


  assign rcache_line[0][140].tag_reg.tag      = reg2hw.tag_140.q;
  assign rcache_line[0][140].tag_reg.qe       = reg2hw.tag_140.qe;
  assign rcache_line[0][140].tag_reg.re       = reg2hw.tag_140.re;
  assign rcache_line[0][140].status_reg.status = reg2hw.status_140.q;//status_reg_t'(reg2hw.status_140.q);
  assign rcache_line[0][140].status_reg.qe    = reg2hw.status_140.qe;
  assign rcache_line[0][140].status_reg.re    = reg2hw.status_140.re;


  assign rcache_line[0][141].tag_reg.tag      = reg2hw.tag_141.q;
  assign rcache_line[0][141].tag_reg.qe       = reg2hw.tag_141.qe;
  assign rcache_line[0][141].tag_reg.re       = reg2hw.tag_141.re;
  assign rcache_line[0][141].status_reg.status = reg2hw.status_141.q;//status_reg_t'(reg2hw.status_141.q);
  assign rcache_line[0][141].status_reg.qe    = reg2hw.status_141.qe;
  assign rcache_line[0][141].status_reg.re    = reg2hw.status_141.re;


  assign rcache_line[0][142].tag_reg.tag      = reg2hw.tag_142.q;
  assign rcache_line[0][142].tag_reg.qe       = reg2hw.tag_142.qe;
  assign rcache_line[0][142].tag_reg.re       = reg2hw.tag_142.re;
  assign rcache_line[0][142].status_reg.status = reg2hw.status_142.q;//status_reg_t'(reg2hw.status_142.q);
  assign rcache_line[0][142].status_reg.qe    = reg2hw.status_142.qe;
  assign rcache_line[0][142].status_reg.re    = reg2hw.status_142.re;


  assign rcache_line[0][143].tag_reg.tag      = reg2hw.tag_143.q;
  assign rcache_line[0][143].tag_reg.qe       = reg2hw.tag_143.qe;
  assign rcache_line[0][143].tag_reg.re       = reg2hw.tag_143.re;
  assign rcache_line[0][143].status_reg.status = reg2hw.status_143.q;//status_reg_t'(reg2hw.status_143.q);
  assign rcache_line[0][143].status_reg.qe    = reg2hw.status_143.qe;
  assign rcache_line[0][143].status_reg.re    = reg2hw.status_143.re;


  assign rcache_line[0][144].tag_reg.tag      = reg2hw.tag_144.q;
  assign rcache_line[0][144].tag_reg.qe       = reg2hw.tag_144.qe;
  assign rcache_line[0][144].tag_reg.re       = reg2hw.tag_144.re;
  assign rcache_line[0][144].status_reg.status = reg2hw.status_144.q;//status_reg_t'(reg2hw.status_144.q);
  assign rcache_line[0][144].status_reg.qe    = reg2hw.status_144.qe;
  assign rcache_line[0][144].status_reg.re    = reg2hw.status_144.re;


  assign rcache_line[0][145].tag_reg.tag      = reg2hw.tag_145.q;
  assign rcache_line[0][145].tag_reg.qe       = reg2hw.tag_145.qe;
  assign rcache_line[0][145].tag_reg.re       = reg2hw.tag_145.re;
  assign rcache_line[0][145].status_reg.status = reg2hw.status_145.q;//status_reg_t'(reg2hw.status_145.q);
  assign rcache_line[0][145].status_reg.qe    = reg2hw.status_145.qe;
  assign rcache_line[0][145].status_reg.re    = reg2hw.status_145.re;


  assign rcache_line[0][146].tag_reg.tag      = reg2hw.tag_146.q;
  assign rcache_line[0][146].tag_reg.qe       = reg2hw.tag_146.qe;
  assign rcache_line[0][146].tag_reg.re       = reg2hw.tag_146.re;
  assign rcache_line[0][146].status_reg.status = reg2hw.status_146.q;//status_reg_t'(reg2hw.status_146.q);
  assign rcache_line[0][146].status_reg.qe    = reg2hw.status_146.qe;
  assign rcache_line[0][146].status_reg.re    = reg2hw.status_146.re;


  assign rcache_line[0][147].tag_reg.tag      = reg2hw.tag_147.q;
  assign rcache_line[0][147].tag_reg.qe       = reg2hw.tag_147.qe;
  assign rcache_line[0][147].tag_reg.re       = reg2hw.tag_147.re;
  assign rcache_line[0][147].status_reg.status = reg2hw.status_147.q;//status_reg_t'(reg2hw.status_147.q);
  assign rcache_line[0][147].status_reg.qe    = reg2hw.status_147.qe;
  assign rcache_line[0][147].status_reg.re    = reg2hw.status_147.re;


  assign rcache_line[0][148].tag_reg.tag      = reg2hw.tag_148.q;
  assign rcache_line[0][148].tag_reg.qe       = reg2hw.tag_148.qe;
  assign rcache_line[0][148].tag_reg.re       = reg2hw.tag_148.re;
  assign rcache_line[0][148].status_reg.status = reg2hw.status_148.q;//status_reg_t'(reg2hw.status_148.q);
  assign rcache_line[0][148].status_reg.qe    = reg2hw.status_148.qe;
  assign rcache_line[0][148].status_reg.re    = reg2hw.status_148.re;


  assign rcache_line[0][149].tag_reg.tag      = reg2hw.tag_149.q;
  assign rcache_line[0][149].tag_reg.qe       = reg2hw.tag_149.qe;
  assign rcache_line[0][149].tag_reg.re       = reg2hw.tag_149.re;
  assign rcache_line[0][149].status_reg.status = reg2hw.status_149.q;//status_reg_t'(reg2hw.status_149.q);
  assign rcache_line[0][149].status_reg.qe    = reg2hw.status_149.qe;
  assign rcache_line[0][149].status_reg.re    = reg2hw.status_149.re;


  assign rcache_line[0][150].tag_reg.tag      = reg2hw.tag_150.q;
  assign rcache_line[0][150].tag_reg.qe       = reg2hw.tag_150.qe;
  assign rcache_line[0][150].tag_reg.re       = reg2hw.tag_150.re;
  assign rcache_line[0][150].status_reg.status = reg2hw.status_150.q;//status_reg_t'(reg2hw.status_150.q);
  assign rcache_line[0][150].status_reg.qe    = reg2hw.status_150.qe;
  assign rcache_line[0][150].status_reg.re    = reg2hw.status_150.re;


  assign rcache_line[0][151].tag_reg.tag      = reg2hw.tag_151.q;
  assign rcache_line[0][151].tag_reg.qe       = reg2hw.tag_151.qe;
  assign rcache_line[0][151].tag_reg.re       = reg2hw.tag_151.re;
  assign rcache_line[0][151].status_reg.status = reg2hw.status_151.q;//status_reg_t'(reg2hw.status_151.q);
  assign rcache_line[0][151].status_reg.qe    = reg2hw.status_151.qe;
  assign rcache_line[0][151].status_reg.re    = reg2hw.status_151.re;


  assign rcache_line[0][152].tag_reg.tag      = reg2hw.tag_152.q;
  assign rcache_line[0][152].tag_reg.qe       = reg2hw.tag_152.qe;
  assign rcache_line[0][152].tag_reg.re       = reg2hw.tag_152.re;
  assign rcache_line[0][152].status_reg.status = reg2hw.status_152.q;//status_reg_t'(reg2hw.status_152.q);
  assign rcache_line[0][152].status_reg.qe    = reg2hw.status_152.qe;
  assign rcache_line[0][152].status_reg.re    = reg2hw.status_152.re;


  assign rcache_line[0][153].tag_reg.tag      = reg2hw.tag_153.q;
  assign rcache_line[0][153].tag_reg.qe       = reg2hw.tag_153.qe;
  assign rcache_line[0][153].tag_reg.re       = reg2hw.tag_153.re;
  assign rcache_line[0][153].status_reg.status = reg2hw.status_153.q;//status_reg_t'(reg2hw.status_153.q);
  assign rcache_line[0][153].status_reg.qe    = reg2hw.status_153.qe;
  assign rcache_line[0][153].status_reg.re    = reg2hw.status_153.re;


  assign rcache_line[0][154].tag_reg.tag      = reg2hw.tag_154.q;
  assign rcache_line[0][154].tag_reg.qe       = reg2hw.tag_154.qe;
  assign rcache_line[0][154].tag_reg.re       = reg2hw.tag_154.re;
  assign rcache_line[0][154].status_reg.status = reg2hw.status_154.q;//status_reg_t'(reg2hw.status_154.q);
  assign rcache_line[0][154].status_reg.qe    = reg2hw.status_154.qe;
  assign rcache_line[0][154].status_reg.re    = reg2hw.status_154.re;


  assign rcache_line[0][155].tag_reg.tag      = reg2hw.tag_155.q;
  assign rcache_line[0][155].tag_reg.qe       = reg2hw.tag_155.qe;
  assign rcache_line[0][155].tag_reg.re       = reg2hw.tag_155.re;
  assign rcache_line[0][155].status_reg.status = reg2hw.status_155.q;//status_reg_t'(reg2hw.status_155.q);
  assign rcache_line[0][155].status_reg.qe    = reg2hw.status_155.qe;
  assign rcache_line[0][155].status_reg.re    = reg2hw.status_155.re;


  assign rcache_line[0][156].tag_reg.tag      = reg2hw.tag_156.q;
  assign rcache_line[0][156].tag_reg.qe       = reg2hw.tag_156.qe;
  assign rcache_line[0][156].tag_reg.re       = reg2hw.tag_156.re;
  assign rcache_line[0][156].status_reg.status = reg2hw.status_156.q;//status_reg_t'(reg2hw.status_156.q);
  assign rcache_line[0][156].status_reg.qe    = reg2hw.status_156.qe;
  assign rcache_line[0][156].status_reg.re    = reg2hw.status_156.re;


  assign rcache_line[0][157].tag_reg.tag      = reg2hw.tag_157.q;
  assign rcache_line[0][157].tag_reg.qe       = reg2hw.tag_157.qe;
  assign rcache_line[0][157].tag_reg.re       = reg2hw.tag_157.re;
  assign rcache_line[0][157].status_reg.status = reg2hw.status_157.q;//status_reg_t'(reg2hw.status_157.q);
  assign rcache_line[0][157].status_reg.qe    = reg2hw.status_157.qe;
  assign rcache_line[0][157].status_reg.re    = reg2hw.status_157.re;


  assign rcache_line[0][158].tag_reg.tag      = reg2hw.tag_158.q;
  assign rcache_line[0][158].tag_reg.qe       = reg2hw.tag_158.qe;
  assign rcache_line[0][158].tag_reg.re       = reg2hw.tag_158.re;
  assign rcache_line[0][158].status_reg.status = reg2hw.status_158.q;//status_reg_t'(reg2hw.status_158.q);
  assign rcache_line[0][158].status_reg.qe    = reg2hw.status_158.qe;
  assign rcache_line[0][158].status_reg.re    = reg2hw.status_158.re;


  assign rcache_line[0][159].tag_reg.tag      = reg2hw.tag_159.q;
  assign rcache_line[0][159].tag_reg.qe       = reg2hw.tag_159.qe;
  assign rcache_line[0][159].tag_reg.re       = reg2hw.tag_159.re;
  assign rcache_line[0][159].status_reg.status = reg2hw.status_159.q;//status_reg_t'(reg2hw.status_159.q);
  assign rcache_line[0][159].status_reg.qe    = reg2hw.status_159.qe;
  assign rcache_line[0][159].status_reg.re    = reg2hw.status_159.re;


  assign rcache_line[0][160].tag_reg.tag      = reg2hw.tag_160.q;
  assign rcache_line[0][160].tag_reg.qe       = reg2hw.tag_160.qe;
  assign rcache_line[0][160].tag_reg.re       = reg2hw.tag_160.re;
  assign rcache_line[0][160].status_reg.status = reg2hw.status_160.q;//status_reg_t'(reg2hw.status_160.q);
  assign rcache_line[0][160].status_reg.qe    = reg2hw.status_160.qe;
  assign rcache_line[0][160].status_reg.re    = reg2hw.status_160.re;


  assign rcache_line[0][161].tag_reg.tag      = reg2hw.tag_161.q;
  assign rcache_line[0][161].tag_reg.qe       = reg2hw.tag_161.qe;
  assign rcache_line[0][161].tag_reg.re       = reg2hw.tag_161.re;
  assign rcache_line[0][161].status_reg.status = reg2hw.status_161.q;//status_reg_t'(reg2hw.status_161.q);
  assign rcache_line[0][161].status_reg.qe    = reg2hw.status_161.qe;
  assign rcache_line[0][161].status_reg.re    = reg2hw.status_161.re;


  assign rcache_line[0][162].tag_reg.tag      = reg2hw.tag_162.q;
  assign rcache_line[0][162].tag_reg.qe       = reg2hw.tag_162.qe;
  assign rcache_line[0][162].tag_reg.re       = reg2hw.tag_162.re;
  assign rcache_line[0][162].status_reg.status = reg2hw.status_162.q;//status_reg_t'(reg2hw.status_162.q);
  assign rcache_line[0][162].status_reg.qe    = reg2hw.status_162.qe;
  assign rcache_line[0][162].status_reg.re    = reg2hw.status_162.re;


  assign rcache_line[0][163].tag_reg.tag      = reg2hw.tag_163.q;
  assign rcache_line[0][163].tag_reg.qe       = reg2hw.tag_163.qe;
  assign rcache_line[0][163].tag_reg.re       = reg2hw.tag_163.re;
  assign rcache_line[0][163].status_reg.status = reg2hw.status_163.q;//status_reg_t'(reg2hw.status_163.q);
  assign rcache_line[0][163].status_reg.qe    = reg2hw.status_163.qe;
  assign rcache_line[0][163].status_reg.re    = reg2hw.status_163.re;


  assign rcache_line[0][164].tag_reg.tag      = reg2hw.tag_164.q;
  assign rcache_line[0][164].tag_reg.qe       = reg2hw.tag_164.qe;
  assign rcache_line[0][164].tag_reg.re       = reg2hw.tag_164.re;
  assign rcache_line[0][164].status_reg.status = reg2hw.status_164.q;//status_reg_t'(reg2hw.status_164.q);
  assign rcache_line[0][164].status_reg.qe    = reg2hw.status_164.qe;
  assign rcache_line[0][164].status_reg.re    = reg2hw.status_164.re;


  assign rcache_line[0][165].tag_reg.tag      = reg2hw.tag_165.q;
  assign rcache_line[0][165].tag_reg.qe       = reg2hw.tag_165.qe;
  assign rcache_line[0][165].tag_reg.re       = reg2hw.tag_165.re;
  assign rcache_line[0][165].status_reg.status = reg2hw.status_165.q;//status_reg_t'(reg2hw.status_165.q);
  assign rcache_line[0][165].status_reg.qe    = reg2hw.status_165.qe;
  assign rcache_line[0][165].status_reg.re    = reg2hw.status_165.re;


  assign rcache_line[0][166].tag_reg.tag      = reg2hw.tag_166.q;
  assign rcache_line[0][166].tag_reg.qe       = reg2hw.tag_166.qe;
  assign rcache_line[0][166].tag_reg.re       = reg2hw.tag_166.re;
  assign rcache_line[0][166].status_reg.status = reg2hw.status_166.q;//status_reg_t'(reg2hw.status_166.q);
  assign rcache_line[0][166].status_reg.qe    = reg2hw.status_166.qe;
  assign rcache_line[0][166].status_reg.re    = reg2hw.status_166.re;


  assign rcache_line[0][167].tag_reg.tag      = reg2hw.tag_167.q;
  assign rcache_line[0][167].tag_reg.qe       = reg2hw.tag_167.qe;
  assign rcache_line[0][167].tag_reg.re       = reg2hw.tag_167.re;
  assign rcache_line[0][167].status_reg.status = reg2hw.status_167.q;//status_reg_t'(reg2hw.status_167.q);
  assign rcache_line[0][167].status_reg.qe    = reg2hw.status_167.qe;
  assign rcache_line[0][167].status_reg.re    = reg2hw.status_167.re;


  assign rcache_line[0][168].tag_reg.tag      = reg2hw.tag_168.q;
  assign rcache_line[0][168].tag_reg.qe       = reg2hw.tag_168.qe;
  assign rcache_line[0][168].tag_reg.re       = reg2hw.tag_168.re;
  assign rcache_line[0][168].status_reg.status = reg2hw.status_168.q;//status_reg_t'(reg2hw.status_168.q);
  assign rcache_line[0][168].status_reg.qe    = reg2hw.status_168.qe;
  assign rcache_line[0][168].status_reg.re    = reg2hw.status_168.re;


  assign rcache_line[0][169].tag_reg.tag      = reg2hw.tag_169.q;
  assign rcache_line[0][169].tag_reg.qe       = reg2hw.tag_169.qe;
  assign rcache_line[0][169].tag_reg.re       = reg2hw.tag_169.re;
  assign rcache_line[0][169].status_reg.status = reg2hw.status_169.q;//status_reg_t'(reg2hw.status_169.q);
  assign rcache_line[0][169].status_reg.qe    = reg2hw.status_169.qe;
  assign rcache_line[0][169].status_reg.re    = reg2hw.status_169.re;


  assign rcache_line[0][170].tag_reg.tag      = reg2hw.tag_170.q;
  assign rcache_line[0][170].tag_reg.qe       = reg2hw.tag_170.qe;
  assign rcache_line[0][170].tag_reg.re       = reg2hw.tag_170.re;
  assign rcache_line[0][170].status_reg.status = reg2hw.status_170.q;//status_reg_t'(reg2hw.status_170.q);
  assign rcache_line[0][170].status_reg.qe    = reg2hw.status_170.qe;
  assign rcache_line[0][170].status_reg.re    = reg2hw.status_170.re;


  assign rcache_line[0][171].tag_reg.tag      = reg2hw.tag_171.q;
  assign rcache_line[0][171].tag_reg.qe       = reg2hw.tag_171.qe;
  assign rcache_line[0][171].tag_reg.re       = reg2hw.tag_171.re;
  assign rcache_line[0][171].status_reg.status = reg2hw.status_171.q;//status_reg_t'(reg2hw.status_171.q);
  assign rcache_line[0][171].status_reg.qe    = reg2hw.status_171.qe;
  assign rcache_line[0][171].status_reg.re    = reg2hw.status_171.re;


  assign rcache_line[0][172].tag_reg.tag      = reg2hw.tag_172.q;
  assign rcache_line[0][172].tag_reg.qe       = reg2hw.tag_172.qe;
  assign rcache_line[0][172].tag_reg.re       = reg2hw.tag_172.re;
  assign rcache_line[0][172].status_reg.status = reg2hw.status_172.q;//status_reg_t'(reg2hw.status_172.q);
  assign rcache_line[0][172].status_reg.qe    = reg2hw.status_172.qe;
  assign rcache_line[0][172].status_reg.re    = reg2hw.status_172.re;


  assign rcache_line[0][173].tag_reg.tag      = reg2hw.tag_173.q;
  assign rcache_line[0][173].tag_reg.qe       = reg2hw.tag_173.qe;
  assign rcache_line[0][173].tag_reg.re       = reg2hw.tag_173.re;
  assign rcache_line[0][173].status_reg.status = reg2hw.status_173.q;//status_reg_t'(reg2hw.status_173.q);
  assign rcache_line[0][173].status_reg.qe    = reg2hw.status_173.qe;
  assign rcache_line[0][173].status_reg.re    = reg2hw.status_173.re;


  assign rcache_line[0][174].tag_reg.tag      = reg2hw.tag_174.q;
  assign rcache_line[0][174].tag_reg.qe       = reg2hw.tag_174.qe;
  assign rcache_line[0][174].tag_reg.re       = reg2hw.tag_174.re;
  assign rcache_line[0][174].status_reg.status = reg2hw.status_174.q;//status_reg_t'(reg2hw.status_174.q);
  assign rcache_line[0][174].status_reg.qe    = reg2hw.status_174.qe;
  assign rcache_line[0][174].status_reg.re    = reg2hw.status_174.re;


  assign rcache_line[0][175].tag_reg.tag      = reg2hw.tag_175.q;
  assign rcache_line[0][175].tag_reg.qe       = reg2hw.tag_175.qe;
  assign rcache_line[0][175].tag_reg.re       = reg2hw.tag_175.re;
  assign rcache_line[0][175].status_reg.status = reg2hw.status_175.q;//status_reg_t'(reg2hw.status_175.q);
  assign rcache_line[0][175].status_reg.qe    = reg2hw.status_175.qe;
  assign rcache_line[0][175].status_reg.re    = reg2hw.status_175.re;


  assign rcache_line[0][176].tag_reg.tag      = reg2hw.tag_176.q;
  assign rcache_line[0][176].tag_reg.qe       = reg2hw.tag_176.qe;
  assign rcache_line[0][176].tag_reg.re       = reg2hw.tag_176.re;
  assign rcache_line[0][176].status_reg.status = reg2hw.status_176.q;//status_reg_t'(reg2hw.status_176.q);
  assign rcache_line[0][176].status_reg.qe    = reg2hw.status_176.qe;
  assign rcache_line[0][176].status_reg.re    = reg2hw.status_176.re;


  assign rcache_line[0][177].tag_reg.tag      = reg2hw.tag_177.q;
  assign rcache_line[0][177].tag_reg.qe       = reg2hw.tag_177.qe;
  assign rcache_line[0][177].tag_reg.re       = reg2hw.tag_177.re;
  assign rcache_line[0][177].status_reg.status = reg2hw.status_177.q;//status_reg_t'(reg2hw.status_177.q);
  assign rcache_line[0][177].status_reg.qe    = reg2hw.status_177.qe;
  assign rcache_line[0][177].status_reg.re    = reg2hw.status_177.re;


  assign rcache_line[0][178].tag_reg.tag      = reg2hw.tag_178.q;
  assign rcache_line[0][178].tag_reg.qe       = reg2hw.tag_178.qe;
  assign rcache_line[0][178].tag_reg.re       = reg2hw.tag_178.re;
  assign rcache_line[0][178].status_reg.status = reg2hw.status_178.q;//status_reg_t'(reg2hw.status_178.q);
  assign rcache_line[0][178].status_reg.qe    = reg2hw.status_178.qe;
  assign rcache_line[0][178].status_reg.re    = reg2hw.status_178.re;


  assign rcache_line[0][179].tag_reg.tag      = reg2hw.tag_179.q;
  assign rcache_line[0][179].tag_reg.qe       = reg2hw.tag_179.qe;
  assign rcache_line[0][179].tag_reg.re       = reg2hw.tag_179.re;
  assign rcache_line[0][179].status_reg.status = reg2hw.status_179.q;//status_reg_t'(reg2hw.status_179.q);
  assign rcache_line[0][179].status_reg.qe    = reg2hw.status_179.qe;
  assign rcache_line[0][179].status_reg.re    = reg2hw.status_179.re;


  assign rcache_line[0][180].tag_reg.tag      = reg2hw.tag_180.q;
  assign rcache_line[0][180].tag_reg.qe       = reg2hw.tag_180.qe;
  assign rcache_line[0][180].tag_reg.re       = reg2hw.tag_180.re;
  assign rcache_line[0][180].status_reg.status = reg2hw.status_180.q;//status_reg_t'(reg2hw.status_180.q);
  assign rcache_line[0][180].status_reg.qe    = reg2hw.status_180.qe;
  assign rcache_line[0][180].status_reg.re    = reg2hw.status_180.re;


  assign rcache_line[0][181].tag_reg.tag      = reg2hw.tag_181.q;
  assign rcache_line[0][181].tag_reg.qe       = reg2hw.tag_181.qe;
  assign rcache_line[0][181].tag_reg.re       = reg2hw.tag_181.re;
  assign rcache_line[0][181].status_reg.status = reg2hw.status_181.q;//status_reg_t'(reg2hw.status_181.q);
  assign rcache_line[0][181].status_reg.qe    = reg2hw.status_181.qe;
  assign rcache_line[0][181].status_reg.re    = reg2hw.status_181.re;


  assign rcache_line[0][182].tag_reg.tag      = reg2hw.tag_182.q;
  assign rcache_line[0][182].tag_reg.qe       = reg2hw.tag_182.qe;
  assign rcache_line[0][182].tag_reg.re       = reg2hw.tag_182.re;
  assign rcache_line[0][182].status_reg.status = reg2hw.status_182.q;//status_reg_t'(reg2hw.status_182.q);
  assign rcache_line[0][182].status_reg.qe    = reg2hw.status_182.qe;
  assign rcache_line[0][182].status_reg.re    = reg2hw.status_182.re;


  assign rcache_line[0][183].tag_reg.tag      = reg2hw.tag_183.q;
  assign rcache_line[0][183].tag_reg.qe       = reg2hw.tag_183.qe;
  assign rcache_line[0][183].tag_reg.re       = reg2hw.tag_183.re;
  assign rcache_line[0][183].status_reg.status = reg2hw.status_183.q;//status_reg_t'(reg2hw.status_183.q);
  assign rcache_line[0][183].status_reg.qe    = reg2hw.status_183.qe;
  assign rcache_line[0][183].status_reg.re    = reg2hw.status_183.re;


  assign rcache_line[0][184].tag_reg.tag      = reg2hw.tag_184.q;
  assign rcache_line[0][184].tag_reg.qe       = reg2hw.tag_184.qe;
  assign rcache_line[0][184].tag_reg.re       = reg2hw.tag_184.re;
  assign rcache_line[0][184].status_reg.status = reg2hw.status_184.q;//status_reg_t'(reg2hw.status_184.q);
  assign rcache_line[0][184].status_reg.qe    = reg2hw.status_184.qe;
  assign rcache_line[0][184].status_reg.re    = reg2hw.status_184.re;


  assign rcache_line[0][185].tag_reg.tag      = reg2hw.tag_185.q;
  assign rcache_line[0][185].tag_reg.qe       = reg2hw.tag_185.qe;
  assign rcache_line[0][185].tag_reg.re       = reg2hw.tag_185.re;
  assign rcache_line[0][185].status_reg.status = reg2hw.status_185.q;//status_reg_t'(reg2hw.status_185.q);
  assign rcache_line[0][185].status_reg.qe    = reg2hw.status_185.qe;
  assign rcache_line[0][185].status_reg.re    = reg2hw.status_185.re;


  assign rcache_line[0][186].tag_reg.tag      = reg2hw.tag_186.q;
  assign rcache_line[0][186].tag_reg.qe       = reg2hw.tag_186.qe;
  assign rcache_line[0][186].tag_reg.re       = reg2hw.tag_186.re;
  assign rcache_line[0][186].status_reg.status = reg2hw.status_186.q;//status_reg_t'(reg2hw.status_186.q);
  assign rcache_line[0][186].status_reg.qe    = reg2hw.status_186.qe;
  assign rcache_line[0][186].status_reg.re    = reg2hw.status_186.re;


  assign rcache_line[0][187].tag_reg.tag      = reg2hw.tag_187.q;
  assign rcache_line[0][187].tag_reg.qe       = reg2hw.tag_187.qe;
  assign rcache_line[0][187].tag_reg.re       = reg2hw.tag_187.re;
  assign rcache_line[0][187].status_reg.status = reg2hw.status_187.q;//status_reg_t'(reg2hw.status_187.q);
  assign rcache_line[0][187].status_reg.qe    = reg2hw.status_187.qe;
  assign rcache_line[0][187].status_reg.re    = reg2hw.status_187.re;


  assign rcache_line[0][188].tag_reg.tag      = reg2hw.tag_188.q;
  assign rcache_line[0][188].tag_reg.qe       = reg2hw.tag_188.qe;
  assign rcache_line[0][188].tag_reg.re       = reg2hw.tag_188.re;
  assign rcache_line[0][188].status_reg.status = reg2hw.status_188.q;//status_reg_t'(reg2hw.status_188.q);
  assign rcache_line[0][188].status_reg.qe    = reg2hw.status_188.qe;
  assign rcache_line[0][188].status_reg.re    = reg2hw.status_188.re;


  assign rcache_line[0][189].tag_reg.tag      = reg2hw.tag_189.q;
  assign rcache_line[0][189].tag_reg.qe       = reg2hw.tag_189.qe;
  assign rcache_line[0][189].tag_reg.re       = reg2hw.tag_189.re;
  assign rcache_line[0][189].status_reg.status = reg2hw.status_189.q;//status_reg_t'(reg2hw.status_189.q);
  assign rcache_line[0][189].status_reg.qe    = reg2hw.status_189.qe;
  assign rcache_line[0][189].status_reg.re    = reg2hw.status_189.re;


  assign rcache_line[0][190].tag_reg.tag      = reg2hw.tag_190.q;
  assign rcache_line[0][190].tag_reg.qe       = reg2hw.tag_190.qe;
  assign rcache_line[0][190].tag_reg.re       = reg2hw.tag_190.re;
  assign rcache_line[0][190].status_reg.status = reg2hw.status_190.q;//status_reg_t'(reg2hw.status_190.q);
  assign rcache_line[0][190].status_reg.qe    = reg2hw.status_190.qe;
  assign rcache_line[0][190].status_reg.re    = reg2hw.status_190.re;


  assign rcache_line[0][191].tag_reg.tag      = reg2hw.tag_191.q;
  assign rcache_line[0][191].tag_reg.qe       = reg2hw.tag_191.qe;
  assign rcache_line[0][191].tag_reg.re       = reg2hw.tag_191.re;
  assign rcache_line[0][191].status_reg.status = reg2hw.status_191.q;//status_reg_t'(reg2hw.status_191.q);
  assign rcache_line[0][191].status_reg.qe    = reg2hw.status_191.qe;
  assign rcache_line[0][191].status_reg.re    = reg2hw.status_191.re;


  assign rcache_line[0][192].tag_reg.tag      = reg2hw.tag_192.q;
  assign rcache_line[0][192].tag_reg.qe       = reg2hw.tag_192.qe;
  assign rcache_line[0][192].tag_reg.re       = reg2hw.tag_192.re;
  assign rcache_line[0][192].status_reg.status = reg2hw.status_192.q;//status_reg_t'(reg2hw.status_192.q);
  assign rcache_line[0][192].status_reg.qe    = reg2hw.status_192.qe;
  assign rcache_line[0][192].status_reg.re    = reg2hw.status_192.re;


  assign rcache_line[0][193].tag_reg.tag      = reg2hw.tag_193.q;
  assign rcache_line[0][193].tag_reg.qe       = reg2hw.tag_193.qe;
  assign rcache_line[0][193].tag_reg.re       = reg2hw.tag_193.re;
  assign rcache_line[0][193].status_reg.status = reg2hw.status_193.q;//status_reg_t'(reg2hw.status_193.q);
  assign rcache_line[0][193].status_reg.qe    = reg2hw.status_193.qe;
  assign rcache_line[0][193].status_reg.re    = reg2hw.status_193.re;


  assign rcache_line[0][194].tag_reg.tag      = reg2hw.tag_194.q;
  assign rcache_line[0][194].tag_reg.qe       = reg2hw.tag_194.qe;
  assign rcache_line[0][194].tag_reg.re       = reg2hw.tag_194.re;
  assign rcache_line[0][194].status_reg.status = reg2hw.status_194.q;//status_reg_t'(reg2hw.status_194.q);
  assign rcache_line[0][194].status_reg.qe    = reg2hw.status_194.qe;
  assign rcache_line[0][194].status_reg.re    = reg2hw.status_194.re;


  assign rcache_line[0][195].tag_reg.tag      = reg2hw.tag_195.q;
  assign rcache_line[0][195].tag_reg.qe       = reg2hw.tag_195.qe;
  assign rcache_line[0][195].tag_reg.re       = reg2hw.tag_195.re;
  assign rcache_line[0][195].status_reg.status = reg2hw.status_195.q;//status_reg_t'(reg2hw.status_195.q);
  assign rcache_line[0][195].status_reg.qe    = reg2hw.status_195.qe;
  assign rcache_line[0][195].status_reg.re    = reg2hw.status_195.re;


  assign rcache_line[0][196].tag_reg.tag      = reg2hw.tag_196.q;
  assign rcache_line[0][196].tag_reg.qe       = reg2hw.tag_196.qe;
  assign rcache_line[0][196].tag_reg.re       = reg2hw.tag_196.re;
  assign rcache_line[0][196].status_reg.status = reg2hw.status_196.q;//status_reg_t'(reg2hw.status_196.q);
  assign rcache_line[0][196].status_reg.qe    = reg2hw.status_196.qe;
  assign rcache_line[0][196].status_reg.re    = reg2hw.status_196.re;


  assign rcache_line[0][197].tag_reg.tag      = reg2hw.tag_197.q;
  assign rcache_line[0][197].tag_reg.qe       = reg2hw.tag_197.qe;
  assign rcache_line[0][197].tag_reg.re       = reg2hw.tag_197.re;
  assign rcache_line[0][197].status_reg.status = reg2hw.status_197.q;//status_reg_t'(reg2hw.status_197.q);
  assign rcache_line[0][197].status_reg.qe    = reg2hw.status_197.qe;
  assign rcache_line[0][197].status_reg.re    = reg2hw.status_197.re;


  assign rcache_line[0][198].tag_reg.tag      = reg2hw.tag_198.q;
  assign rcache_line[0][198].tag_reg.qe       = reg2hw.tag_198.qe;
  assign rcache_line[0][198].tag_reg.re       = reg2hw.tag_198.re;
  assign rcache_line[0][198].status_reg.status = reg2hw.status_198.q;//status_reg_t'(reg2hw.status_198.q);
  assign rcache_line[0][198].status_reg.qe    = reg2hw.status_198.qe;
  assign rcache_line[0][198].status_reg.re    = reg2hw.status_198.re;


  assign rcache_line[0][199].tag_reg.tag      = reg2hw.tag_199.q;
  assign rcache_line[0][199].tag_reg.qe       = reg2hw.tag_199.qe;
  assign rcache_line[0][199].tag_reg.re       = reg2hw.tag_199.re;
  assign rcache_line[0][199].status_reg.status = reg2hw.status_199.q;//status_reg_t'(reg2hw.status_199.q);
  assign rcache_line[0][199].status_reg.qe    = reg2hw.status_199.qe;
  assign rcache_line[0][199].status_reg.re    = reg2hw.status_199.re;


  assign rcache_line[0][200].tag_reg.tag      = reg2hw.tag_200.q;
  assign rcache_line[0][200].tag_reg.qe       = reg2hw.tag_200.qe;
  assign rcache_line[0][200].tag_reg.re       = reg2hw.tag_200.re;
  assign rcache_line[0][200].status_reg.status = reg2hw.status_200.q;//status_reg_t'(reg2hw.status_200.q);
  assign rcache_line[0][200].status_reg.qe    = reg2hw.status_200.qe;
  assign rcache_line[0][200].status_reg.re    = reg2hw.status_200.re;


  assign rcache_line[0][201].tag_reg.tag      = reg2hw.tag_201.q;
  assign rcache_line[0][201].tag_reg.qe       = reg2hw.tag_201.qe;
  assign rcache_line[0][201].tag_reg.re       = reg2hw.tag_201.re;
  assign rcache_line[0][201].status_reg.status = reg2hw.status_201.q;//status_reg_t'(reg2hw.status_201.q);
  assign rcache_line[0][201].status_reg.qe    = reg2hw.status_201.qe;
  assign rcache_line[0][201].status_reg.re    = reg2hw.status_201.re;


  assign rcache_line[0][202].tag_reg.tag      = reg2hw.tag_202.q;
  assign rcache_line[0][202].tag_reg.qe       = reg2hw.tag_202.qe;
  assign rcache_line[0][202].tag_reg.re       = reg2hw.tag_202.re;
  assign rcache_line[0][202].status_reg.status = reg2hw.status_202.q;//status_reg_t'(reg2hw.status_202.q);
  assign rcache_line[0][202].status_reg.qe    = reg2hw.status_202.qe;
  assign rcache_line[0][202].status_reg.re    = reg2hw.status_202.re;


  assign rcache_line[0][203].tag_reg.tag      = reg2hw.tag_203.q;
  assign rcache_line[0][203].tag_reg.qe       = reg2hw.tag_203.qe;
  assign rcache_line[0][203].tag_reg.re       = reg2hw.tag_203.re;
  assign rcache_line[0][203].status_reg.status = reg2hw.status_203.q;//status_reg_t'(reg2hw.status_203.q);
  assign rcache_line[0][203].status_reg.qe    = reg2hw.status_203.qe;
  assign rcache_line[0][203].status_reg.re    = reg2hw.status_203.re;


  assign rcache_line[0][204].tag_reg.tag      = reg2hw.tag_204.q;
  assign rcache_line[0][204].tag_reg.qe       = reg2hw.tag_204.qe;
  assign rcache_line[0][204].tag_reg.re       = reg2hw.tag_204.re;
  assign rcache_line[0][204].status_reg.status = reg2hw.status_204.q;//status_reg_t'(reg2hw.status_204.q);
  assign rcache_line[0][204].status_reg.qe    = reg2hw.status_204.qe;
  assign rcache_line[0][204].status_reg.re    = reg2hw.status_204.re;


  assign rcache_line[0][205].tag_reg.tag      = reg2hw.tag_205.q;
  assign rcache_line[0][205].tag_reg.qe       = reg2hw.tag_205.qe;
  assign rcache_line[0][205].tag_reg.re       = reg2hw.tag_205.re;
  assign rcache_line[0][205].status_reg.status = reg2hw.status_205.q;//status_reg_t'(reg2hw.status_205.q);
  assign rcache_line[0][205].status_reg.qe    = reg2hw.status_205.qe;
  assign rcache_line[0][205].status_reg.re    = reg2hw.status_205.re;


  assign rcache_line[0][206].tag_reg.tag      = reg2hw.tag_206.q;
  assign rcache_line[0][206].tag_reg.qe       = reg2hw.tag_206.qe;
  assign rcache_line[0][206].tag_reg.re       = reg2hw.tag_206.re;
  assign rcache_line[0][206].status_reg.status = reg2hw.status_206.q;//status_reg_t'(reg2hw.status_206.q);
  assign rcache_line[0][206].status_reg.qe    = reg2hw.status_206.qe;
  assign rcache_line[0][206].status_reg.re    = reg2hw.status_206.re;


  assign rcache_line[0][207].tag_reg.tag      = reg2hw.tag_207.q;
  assign rcache_line[0][207].tag_reg.qe       = reg2hw.tag_207.qe;
  assign rcache_line[0][207].tag_reg.re       = reg2hw.tag_207.re;
  assign rcache_line[0][207].status_reg.status = reg2hw.status_207.q;//status_reg_t'(reg2hw.status_207.q);
  assign rcache_line[0][207].status_reg.qe    = reg2hw.status_207.qe;
  assign rcache_line[0][207].status_reg.re    = reg2hw.status_207.re;


  assign rcache_line[0][208].tag_reg.tag      = reg2hw.tag_208.q;
  assign rcache_line[0][208].tag_reg.qe       = reg2hw.tag_208.qe;
  assign rcache_line[0][208].tag_reg.re       = reg2hw.tag_208.re;
  assign rcache_line[0][208].status_reg.status = reg2hw.status_208.q;//status_reg_t'(reg2hw.status_208.q);
  assign rcache_line[0][208].status_reg.qe    = reg2hw.status_208.qe;
  assign rcache_line[0][208].status_reg.re    = reg2hw.status_208.re;


  assign rcache_line[0][209].tag_reg.tag      = reg2hw.tag_209.q;
  assign rcache_line[0][209].tag_reg.qe       = reg2hw.tag_209.qe;
  assign rcache_line[0][209].tag_reg.re       = reg2hw.tag_209.re;
  assign rcache_line[0][209].status_reg.status = reg2hw.status_209.q;//status_reg_t'(reg2hw.status_209.q);
  assign rcache_line[0][209].status_reg.qe    = reg2hw.status_209.qe;
  assign rcache_line[0][209].status_reg.re    = reg2hw.status_209.re;


  assign rcache_line[0][210].tag_reg.tag      = reg2hw.tag_210.q;
  assign rcache_line[0][210].tag_reg.qe       = reg2hw.tag_210.qe;
  assign rcache_line[0][210].tag_reg.re       = reg2hw.tag_210.re;
  assign rcache_line[0][210].status_reg.status = reg2hw.status_210.q;//status_reg_t'(reg2hw.status_210.q);
  assign rcache_line[0][210].status_reg.qe    = reg2hw.status_210.qe;
  assign rcache_line[0][210].status_reg.re    = reg2hw.status_210.re;


  assign rcache_line[0][211].tag_reg.tag      = reg2hw.tag_211.q;
  assign rcache_line[0][211].tag_reg.qe       = reg2hw.tag_211.qe;
  assign rcache_line[0][211].tag_reg.re       = reg2hw.tag_211.re;
  assign rcache_line[0][211].status_reg.status = reg2hw.status_211.q;//status_reg_t'(reg2hw.status_211.q);
  assign rcache_line[0][211].status_reg.qe    = reg2hw.status_211.qe;
  assign rcache_line[0][211].status_reg.re    = reg2hw.status_211.re;


  assign rcache_line[0][212].tag_reg.tag      = reg2hw.tag_212.q;
  assign rcache_line[0][212].tag_reg.qe       = reg2hw.tag_212.qe;
  assign rcache_line[0][212].tag_reg.re       = reg2hw.tag_212.re;
  assign rcache_line[0][212].status_reg.status = reg2hw.status_212.q;//status_reg_t'(reg2hw.status_212.q);
  assign rcache_line[0][212].status_reg.qe    = reg2hw.status_212.qe;
  assign rcache_line[0][212].status_reg.re    = reg2hw.status_212.re;


  assign rcache_line[0][213].tag_reg.tag      = reg2hw.tag_213.q;
  assign rcache_line[0][213].tag_reg.qe       = reg2hw.tag_213.qe;
  assign rcache_line[0][213].tag_reg.re       = reg2hw.tag_213.re;
  assign rcache_line[0][213].status_reg.status = reg2hw.status_213.q;//status_reg_t'(reg2hw.status_213.q);
  assign rcache_line[0][213].status_reg.qe    = reg2hw.status_213.qe;
  assign rcache_line[0][213].status_reg.re    = reg2hw.status_213.re;


  assign rcache_line[0][214].tag_reg.tag      = reg2hw.tag_214.q;
  assign rcache_line[0][214].tag_reg.qe       = reg2hw.tag_214.qe;
  assign rcache_line[0][214].tag_reg.re       = reg2hw.tag_214.re;
  assign rcache_line[0][214].status_reg.status = reg2hw.status_214.q;//status_reg_t'(reg2hw.status_214.q);
  assign rcache_line[0][214].status_reg.qe    = reg2hw.status_214.qe;
  assign rcache_line[0][214].status_reg.re    = reg2hw.status_214.re;


  assign rcache_line[0][215].tag_reg.tag      = reg2hw.tag_215.q;
  assign rcache_line[0][215].tag_reg.qe       = reg2hw.tag_215.qe;
  assign rcache_line[0][215].tag_reg.re       = reg2hw.tag_215.re;
  assign rcache_line[0][215].status_reg.status = reg2hw.status_215.q;//status_reg_t'(reg2hw.status_215.q);
  assign rcache_line[0][215].status_reg.qe    = reg2hw.status_215.qe;
  assign rcache_line[0][215].status_reg.re    = reg2hw.status_215.re;


  assign rcache_line[0][216].tag_reg.tag      = reg2hw.tag_216.q;
  assign rcache_line[0][216].tag_reg.qe       = reg2hw.tag_216.qe;
  assign rcache_line[0][216].tag_reg.re       = reg2hw.tag_216.re;
  assign rcache_line[0][216].status_reg.status = reg2hw.status_216.q;//status_reg_t'(reg2hw.status_216.q);
  assign rcache_line[0][216].status_reg.qe    = reg2hw.status_216.qe;
  assign rcache_line[0][216].status_reg.re    = reg2hw.status_216.re;


  assign rcache_line[0][217].tag_reg.tag      = reg2hw.tag_217.q;
  assign rcache_line[0][217].tag_reg.qe       = reg2hw.tag_217.qe;
  assign rcache_line[0][217].tag_reg.re       = reg2hw.tag_217.re;
  assign rcache_line[0][217].status_reg.status = reg2hw.status_217.q;//status_reg_t'(reg2hw.status_217.q);
  assign rcache_line[0][217].status_reg.qe    = reg2hw.status_217.qe;
  assign rcache_line[0][217].status_reg.re    = reg2hw.status_217.re;


  assign rcache_line[0][218].tag_reg.tag      = reg2hw.tag_218.q;
  assign rcache_line[0][218].tag_reg.qe       = reg2hw.tag_218.qe;
  assign rcache_line[0][218].tag_reg.re       = reg2hw.tag_218.re;
  assign rcache_line[0][218].status_reg.status = reg2hw.status_218.q;//status_reg_t'(reg2hw.status_218.q);
  assign rcache_line[0][218].status_reg.qe    = reg2hw.status_218.qe;
  assign rcache_line[0][218].status_reg.re    = reg2hw.status_218.re;


  assign rcache_line[0][219].tag_reg.tag      = reg2hw.tag_219.q;
  assign rcache_line[0][219].tag_reg.qe       = reg2hw.tag_219.qe;
  assign rcache_line[0][219].tag_reg.re       = reg2hw.tag_219.re;
  assign rcache_line[0][219].status_reg.status = reg2hw.status_219.q;//status_reg_t'(reg2hw.status_219.q);
  assign rcache_line[0][219].status_reg.qe    = reg2hw.status_219.qe;
  assign rcache_line[0][219].status_reg.re    = reg2hw.status_219.re;


  assign rcache_line[0][220].tag_reg.tag      = reg2hw.tag_220.q;
  assign rcache_line[0][220].tag_reg.qe       = reg2hw.tag_220.qe;
  assign rcache_line[0][220].tag_reg.re       = reg2hw.tag_220.re;
  assign rcache_line[0][220].status_reg.status = reg2hw.status_220.q;//status_reg_t'(reg2hw.status_220.q);
  assign rcache_line[0][220].status_reg.qe    = reg2hw.status_220.qe;
  assign rcache_line[0][220].status_reg.re    = reg2hw.status_220.re;


  assign rcache_line[0][221].tag_reg.tag      = reg2hw.tag_221.q;
  assign rcache_line[0][221].tag_reg.qe       = reg2hw.tag_221.qe;
  assign rcache_line[0][221].tag_reg.re       = reg2hw.tag_221.re;
  assign rcache_line[0][221].status_reg.status = reg2hw.status_221.q;//status_reg_t'(reg2hw.status_221.q);
  assign rcache_line[0][221].status_reg.qe    = reg2hw.status_221.qe;
  assign rcache_line[0][221].status_reg.re    = reg2hw.status_221.re;


  assign rcache_line[0][222].tag_reg.tag      = reg2hw.tag_222.q;
  assign rcache_line[0][222].tag_reg.qe       = reg2hw.tag_222.qe;
  assign rcache_line[0][222].tag_reg.re       = reg2hw.tag_222.re;
  assign rcache_line[0][222].status_reg.status = reg2hw.status_222.q;//status_reg_t'(reg2hw.status_222.q);
  assign rcache_line[0][222].status_reg.qe    = reg2hw.status_222.qe;
  assign rcache_line[0][222].status_reg.re    = reg2hw.status_222.re;


  assign rcache_line[0][223].tag_reg.tag      = reg2hw.tag_223.q;
  assign rcache_line[0][223].tag_reg.qe       = reg2hw.tag_223.qe;
  assign rcache_line[0][223].tag_reg.re       = reg2hw.tag_223.re;
  assign rcache_line[0][223].status_reg.status = reg2hw.status_223.q;//status_reg_t'(reg2hw.status_223.q);
  assign rcache_line[0][223].status_reg.qe    = reg2hw.status_223.qe;
  assign rcache_line[0][223].status_reg.re    = reg2hw.status_223.re;


  assign rcache_line[0][224].tag_reg.tag      = reg2hw.tag_224.q;
  assign rcache_line[0][224].tag_reg.qe       = reg2hw.tag_224.qe;
  assign rcache_line[0][224].tag_reg.re       = reg2hw.tag_224.re;
  assign rcache_line[0][224].status_reg.status = reg2hw.status_224.q;//status_reg_t'(reg2hw.status_224.q);
  assign rcache_line[0][224].status_reg.qe    = reg2hw.status_224.qe;
  assign rcache_line[0][224].status_reg.re    = reg2hw.status_224.re;


  assign rcache_line[0][225].tag_reg.tag      = reg2hw.tag_225.q;
  assign rcache_line[0][225].tag_reg.qe       = reg2hw.tag_225.qe;
  assign rcache_line[0][225].tag_reg.re       = reg2hw.tag_225.re;
  assign rcache_line[0][225].status_reg.status = reg2hw.status_225.q;//status_reg_t'(reg2hw.status_225.q);
  assign rcache_line[0][225].status_reg.qe    = reg2hw.status_225.qe;
  assign rcache_line[0][225].status_reg.re    = reg2hw.status_225.re;


  assign rcache_line[0][226].tag_reg.tag      = reg2hw.tag_226.q;
  assign rcache_line[0][226].tag_reg.qe       = reg2hw.tag_226.qe;
  assign rcache_line[0][226].tag_reg.re       = reg2hw.tag_226.re;
  assign rcache_line[0][226].status_reg.status = reg2hw.status_226.q;//status_reg_t'(reg2hw.status_226.q);
  assign rcache_line[0][226].status_reg.qe    = reg2hw.status_226.qe;
  assign rcache_line[0][226].status_reg.re    = reg2hw.status_226.re;


  assign rcache_line[0][227].tag_reg.tag      = reg2hw.tag_227.q;
  assign rcache_line[0][227].tag_reg.qe       = reg2hw.tag_227.qe;
  assign rcache_line[0][227].tag_reg.re       = reg2hw.tag_227.re;
  assign rcache_line[0][227].status_reg.status = reg2hw.status_227.q;//status_reg_t'(reg2hw.status_227.q);
  assign rcache_line[0][227].status_reg.qe    = reg2hw.status_227.qe;
  assign rcache_line[0][227].status_reg.re    = reg2hw.status_227.re;


  assign rcache_line[0][228].tag_reg.tag      = reg2hw.tag_228.q;
  assign rcache_line[0][228].tag_reg.qe       = reg2hw.tag_228.qe;
  assign rcache_line[0][228].tag_reg.re       = reg2hw.tag_228.re;
  assign rcache_line[0][228].status_reg.status = reg2hw.status_228.q;//status_reg_t'(reg2hw.status_228.q);
  assign rcache_line[0][228].status_reg.qe    = reg2hw.status_228.qe;
  assign rcache_line[0][228].status_reg.re    = reg2hw.status_228.re;


  assign rcache_line[0][229].tag_reg.tag      = reg2hw.tag_229.q;
  assign rcache_line[0][229].tag_reg.qe       = reg2hw.tag_229.qe;
  assign rcache_line[0][229].tag_reg.re       = reg2hw.tag_229.re;
  assign rcache_line[0][229].status_reg.status = reg2hw.status_229.q;//status_reg_t'(reg2hw.status_229.q);
  assign rcache_line[0][229].status_reg.qe    = reg2hw.status_229.qe;
  assign rcache_line[0][229].status_reg.re    = reg2hw.status_229.re;


  assign rcache_line[0][230].tag_reg.tag      = reg2hw.tag_230.q;
  assign rcache_line[0][230].tag_reg.qe       = reg2hw.tag_230.qe;
  assign rcache_line[0][230].tag_reg.re       = reg2hw.tag_230.re;
  assign rcache_line[0][230].status_reg.status = reg2hw.status_230.q;//status_reg_t'(reg2hw.status_230.q);
  assign rcache_line[0][230].status_reg.qe    = reg2hw.status_230.qe;
  assign rcache_line[0][230].status_reg.re    = reg2hw.status_230.re;


  assign rcache_line[0][231].tag_reg.tag      = reg2hw.tag_231.q;
  assign rcache_line[0][231].tag_reg.qe       = reg2hw.tag_231.qe;
  assign rcache_line[0][231].tag_reg.re       = reg2hw.tag_231.re;
  assign rcache_line[0][231].status_reg.status = reg2hw.status_231.q;//status_reg_t'(reg2hw.status_231.q);
  assign rcache_line[0][231].status_reg.qe    = reg2hw.status_231.qe;
  assign rcache_line[0][231].status_reg.re    = reg2hw.status_231.re;


  assign rcache_line[0][232].tag_reg.tag      = reg2hw.tag_232.q;
  assign rcache_line[0][232].tag_reg.qe       = reg2hw.tag_232.qe;
  assign rcache_line[0][232].tag_reg.re       = reg2hw.tag_232.re;
  assign rcache_line[0][232].status_reg.status = reg2hw.status_232.q;//status_reg_t'(reg2hw.status_232.q);
  assign rcache_line[0][232].status_reg.qe    = reg2hw.status_232.qe;
  assign rcache_line[0][232].status_reg.re    = reg2hw.status_232.re;


  assign rcache_line[0][233].tag_reg.tag      = reg2hw.tag_233.q;
  assign rcache_line[0][233].tag_reg.qe       = reg2hw.tag_233.qe;
  assign rcache_line[0][233].tag_reg.re       = reg2hw.tag_233.re;
  assign rcache_line[0][233].status_reg.status = reg2hw.status_233.q;//status_reg_t'(reg2hw.status_233.q);
  assign rcache_line[0][233].status_reg.qe    = reg2hw.status_233.qe;
  assign rcache_line[0][233].status_reg.re    = reg2hw.status_233.re;


  assign rcache_line[0][234].tag_reg.tag      = reg2hw.tag_234.q;
  assign rcache_line[0][234].tag_reg.qe       = reg2hw.tag_234.qe;
  assign rcache_line[0][234].tag_reg.re       = reg2hw.tag_234.re;
  assign rcache_line[0][234].status_reg.status = reg2hw.status_234.q;//status_reg_t'(reg2hw.status_234.q);
  assign rcache_line[0][234].status_reg.qe    = reg2hw.status_234.qe;
  assign rcache_line[0][234].status_reg.re    = reg2hw.status_234.re;


  assign rcache_line[0][235].tag_reg.tag      = reg2hw.tag_235.q;
  assign rcache_line[0][235].tag_reg.qe       = reg2hw.tag_235.qe;
  assign rcache_line[0][235].tag_reg.re       = reg2hw.tag_235.re;
  assign rcache_line[0][235].status_reg.status = reg2hw.status_235.q;//status_reg_t'(reg2hw.status_235.q);
  assign rcache_line[0][235].status_reg.qe    = reg2hw.status_235.qe;
  assign rcache_line[0][235].status_reg.re    = reg2hw.status_235.re;


  assign rcache_line[0][236].tag_reg.tag      = reg2hw.tag_236.q;
  assign rcache_line[0][236].tag_reg.qe       = reg2hw.tag_236.qe;
  assign rcache_line[0][236].tag_reg.re       = reg2hw.tag_236.re;
  assign rcache_line[0][236].status_reg.status = reg2hw.status_236.q;//status_reg_t'(reg2hw.status_236.q);
  assign rcache_line[0][236].status_reg.qe    = reg2hw.status_236.qe;
  assign rcache_line[0][236].status_reg.re    = reg2hw.status_236.re;


  assign rcache_line[0][237].tag_reg.tag      = reg2hw.tag_237.q;
  assign rcache_line[0][237].tag_reg.qe       = reg2hw.tag_237.qe;
  assign rcache_line[0][237].tag_reg.re       = reg2hw.tag_237.re;
  assign rcache_line[0][237].status_reg.status = reg2hw.status_237.q;//status_reg_t'(reg2hw.status_237.q);
  assign rcache_line[0][237].status_reg.qe    = reg2hw.status_237.qe;
  assign rcache_line[0][237].status_reg.re    = reg2hw.status_237.re;


  assign rcache_line[0][238].tag_reg.tag      = reg2hw.tag_238.q;
  assign rcache_line[0][238].tag_reg.qe       = reg2hw.tag_238.qe;
  assign rcache_line[0][238].tag_reg.re       = reg2hw.tag_238.re;
  assign rcache_line[0][238].status_reg.status = reg2hw.status_238.q;//status_reg_t'(reg2hw.status_238.q);
  assign rcache_line[0][238].status_reg.qe    = reg2hw.status_238.qe;
  assign rcache_line[0][238].status_reg.re    = reg2hw.status_238.re;


  assign rcache_line[0][239].tag_reg.tag      = reg2hw.tag_239.q;
  assign rcache_line[0][239].tag_reg.qe       = reg2hw.tag_239.qe;
  assign rcache_line[0][239].tag_reg.re       = reg2hw.tag_239.re;
  assign rcache_line[0][239].status_reg.status = reg2hw.status_239.q;//status_reg_t'(reg2hw.status_239.q);
  assign rcache_line[0][239].status_reg.qe    = reg2hw.status_239.qe;
  assign rcache_line[0][239].status_reg.re    = reg2hw.status_239.re;


  assign rcache_line[0][240].tag_reg.tag      = reg2hw.tag_240.q;
  assign rcache_line[0][240].tag_reg.qe       = reg2hw.tag_240.qe;
  assign rcache_line[0][240].tag_reg.re       = reg2hw.tag_240.re;
  assign rcache_line[0][240].status_reg.status = reg2hw.status_240.q;//status_reg_t'(reg2hw.status_240.q);
  assign rcache_line[0][240].status_reg.qe    = reg2hw.status_240.qe;
  assign rcache_line[0][240].status_reg.re    = reg2hw.status_240.re;


  assign rcache_line[0][241].tag_reg.tag      = reg2hw.tag_241.q;
  assign rcache_line[0][241].tag_reg.qe       = reg2hw.tag_241.qe;
  assign rcache_line[0][241].tag_reg.re       = reg2hw.tag_241.re;
  assign rcache_line[0][241].status_reg.status = reg2hw.status_241.q;//status_reg_t'(reg2hw.status_241.q);
  assign rcache_line[0][241].status_reg.qe    = reg2hw.status_241.qe;
  assign rcache_line[0][241].status_reg.re    = reg2hw.status_241.re;


  assign rcache_line[0][242].tag_reg.tag      = reg2hw.tag_242.q;
  assign rcache_line[0][242].tag_reg.qe       = reg2hw.tag_242.qe;
  assign rcache_line[0][242].tag_reg.re       = reg2hw.tag_242.re;
  assign rcache_line[0][242].status_reg.status = reg2hw.status_242.q;//status_reg_t'(reg2hw.status_242.q);
  assign rcache_line[0][242].status_reg.qe    = reg2hw.status_242.qe;
  assign rcache_line[0][242].status_reg.re    = reg2hw.status_242.re;


  assign rcache_line[0][243].tag_reg.tag      = reg2hw.tag_243.q;
  assign rcache_line[0][243].tag_reg.qe       = reg2hw.tag_243.qe;
  assign rcache_line[0][243].tag_reg.re       = reg2hw.tag_243.re;
  assign rcache_line[0][243].status_reg.status = reg2hw.status_243.q;//status_reg_t'(reg2hw.status_243.q);
  assign rcache_line[0][243].status_reg.qe    = reg2hw.status_243.qe;
  assign rcache_line[0][243].status_reg.re    = reg2hw.status_243.re;


  assign rcache_line[0][244].tag_reg.tag      = reg2hw.tag_244.q;
  assign rcache_line[0][244].tag_reg.qe       = reg2hw.tag_244.qe;
  assign rcache_line[0][244].tag_reg.re       = reg2hw.tag_244.re;
  assign rcache_line[0][244].status_reg.status = reg2hw.status_244.q;//status_reg_t'(reg2hw.status_244.q);
  assign rcache_line[0][244].status_reg.qe    = reg2hw.status_244.qe;
  assign rcache_line[0][244].status_reg.re    = reg2hw.status_244.re;


  assign rcache_line[0][245].tag_reg.tag      = reg2hw.tag_245.q;
  assign rcache_line[0][245].tag_reg.qe       = reg2hw.tag_245.qe;
  assign rcache_line[0][245].tag_reg.re       = reg2hw.tag_245.re;
  assign rcache_line[0][245].status_reg.status = reg2hw.status_245.q;//status_reg_t'(reg2hw.status_245.q);
  assign rcache_line[0][245].status_reg.qe    = reg2hw.status_245.qe;
  assign rcache_line[0][245].status_reg.re    = reg2hw.status_245.re;


  assign rcache_line[0][246].tag_reg.tag      = reg2hw.tag_246.q;
  assign rcache_line[0][246].tag_reg.qe       = reg2hw.tag_246.qe;
  assign rcache_line[0][246].tag_reg.re       = reg2hw.tag_246.re;
  assign rcache_line[0][246].status_reg.status = reg2hw.status_246.q;//status_reg_t'(reg2hw.status_246.q);
  assign rcache_line[0][246].status_reg.qe    = reg2hw.status_246.qe;
  assign rcache_line[0][246].status_reg.re    = reg2hw.status_246.re;


  assign rcache_line[0][247].tag_reg.tag      = reg2hw.tag_247.q;
  assign rcache_line[0][247].tag_reg.qe       = reg2hw.tag_247.qe;
  assign rcache_line[0][247].tag_reg.re       = reg2hw.tag_247.re;
  assign rcache_line[0][247].status_reg.status = reg2hw.status_247.q;//status_reg_t'(reg2hw.status_247.q);
  assign rcache_line[0][247].status_reg.qe    = reg2hw.status_247.qe;
  assign rcache_line[0][247].status_reg.re    = reg2hw.status_247.re;


  assign rcache_line[0][248].tag_reg.tag      = reg2hw.tag_248.q;
  assign rcache_line[0][248].tag_reg.qe       = reg2hw.tag_248.qe;
  assign rcache_line[0][248].tag_reg.re       = reg2hw.tag_248.re;
  assign rcache_line[0][248].status_reg.status = reg2hw.status_248.q;//status_reg_t'(reg2hw.status_248.q);
  assign rcache_line[0][248].status_reg.qe    = reg2hw.status_248.qe;
  assign rcache_line[0][248].status_reg.re    = reg2hw.status_248.re;


  assign rcache_line[0][249].tag_reg.tag      = reg2hw.tag_249.q;
  assign rcache_line[0][249].tag_reg.qe       = reg2hw.tag_249.qe;
  assign rcache_line[0][249].tag_reg.re       = reg2hw.tag_249.re;
  assign rcache_line[0][249].status_reg.status = reg2hw.status_249.q;//status_reg_t'(reg2hw.status_249.q);
  assign rcache_line[0][249].status_reg.qe    = reg2hw.status_249.qe;
  assign rcache_line[0][249].status_reg.re    = reg2hw.status_249.re;


  assign rcache_line[0][250].tag_reg.tag      = reg2hw.tag_250.q;
  assign rcache_line[0][250].tag_reg.qe       = reg2hw.tag_250.qe;
  assign rcache_line[0][250].tag_reg.re       = reg2hw.tag_250.re;
  assign rcache_line[0][250].status_reg.status = reg2hw.status_250.q;//status_reg_t'(reg2hw.status_250.q);
  assign rcache_line[0][250].status_reg.qe    = reg2hw.status_250.qe;
  assign rcache_line[0][250].status_reg.re    = reg2hw.status_250.re;


  assign rcache_line[0][251].tag_reg.tag      = reg2hw.tag_251.q;
  assign rcache_line[0][251].tag_reg.qe       = reg2hw.tag_251.qe;
  assign rcache_line[0][251].tag_reg.re       = reg2hw.tag_251.re;
  assign rcache_line[0][251].status_reg.status = reg2hw.status_251.q;//status_reg_t'(reg2hw.status_251.q);
  assign rcache_line[0][251].status_reg.qe    = reg2hw.status_251.qe;
  assign rcache_line[0][251].status_reg.re    = reg2hw.status_251.re;


  assign rcache_line[0][252].tag_reg.tag      = reg2hw.tag_252.q;
  assign rcache_line[0][252].tag_reg.qe       = reg2hw.tag_252.qe;
  assign rcache_line[0][252].tag_reg.re       = reg2hw.tag_252.re;
  assign rcache_line[0][252].status_reg.status = reg2hw.status_252.q;//status_reg_t'(reg2hw.status_252.q);
  assign rcache_line[0][252].status_reg.qe    = reg2hw.status_252.qe;
  assign rcache_line[0][252].status_reg.re    = reg2hw.status_252.re;


  assign rcache_line[0][253].tag_reg.tag      = reg2hw.tag_253.q;
  assign rcache_line[0][253].tag_reg.qe       = reg2hw.tag_253.qe;
  assign rcache_line[0][253].tag_reg.re       = reg2hw.tag_253.re;
  assign rcache_line[0][253].status_reg.status = reg2hw.status_253.q;//status_reg_t'(reg2hw.status_253.q);
  assign rcache_line[0][253].status_reg.qe    = reg2hw.status_253.qe;
  assign rcache_line[0][253].status_reg.re    = reg2hw.status_253.re;


  assign rcache_line[0][254].tag_reg.tag      = reg2hw.tag_254.q;
  assign rcache_line[0][254].tag_reg.qe       = reg2hw.tag_254.qe;
  assign rcache_line[0][254].tag_reg.re       = reg2hw.tag_254.re;
  assign rcache_line[0][254].status_reg.status = reg2hw.status_254.q;//status_reg_t'(reg2hw.status_254.q);
  assign rcache_line[0][254].status_reg.qe    = reg2hw.status_254.qe;
  assign rcache_line[0][254].status_reg.re    = reg2hw.status_254.re;


  assign rcache_line[0][255].tag_reg.tag      = reg2hw.tag_255.q;
  assign rcache_line[0][255].tag_reg.qe       = reg2hw.tag_255.qe;
  assign rcache_line[0][255].tag_reg.re       = reg2hw.tag_255.re;
  assign rcache_line[0][255].status_reg.status = reg2hw.status_255.q;//status_reg_t'(reg2hw.status_255.q);
  assign rcache_line[0][255].status_reg.qe    = reg2hw.status_255.qe;
  assign rcache_line[0][255].status_reg.re    = reg2hw.status_255.re;


  assign rcache_line[1][0].tag_reg.tag      = reg2hw.tag_256.q;
  assign rcache_line[1][0].tag_reg.qe       = reg2hw.tag_256.qe;
  assign rcache_line[1][0].tag_reg.re       = reg2hw.tag_256.re;
  assign rcache_line[1][0].status_reg.status = reg2hw.status_256.q;//status_reg_t'(reg2hw.status_256.q);
  assign rcache_line[1][0].status_reg.qe    = reg2hw.status_256.qe;
  assign rcache_line[1][0].status_reg.re    = reg2hw.status_256.re;


  assign rcache_line[1][1].tag_reg.tag      = reg2hw.tag_257.q;
  assign rcache_line[1][1].tag_reg.qe       = reg2hw.tag_257.qe;
  assign rcache_line[1][1].tag_reg.re       = reg2hw.tag_257.re;
  assign rcache_line[1][1].status_reg.status = reg2hw.status_257.q;//status_reg_t'(reg2hw.status_257.q);
  assign rcache_line[1][1].status_reg.qe    = reg2hw.status_257.qe;
  assign rcache_line[1][1].status_reg.re    = reg2hw.status_257.re;


  assign rcache_line[1][2].tag_reg.tag      = reg2hw.tag_258.q;
  assign rcache_line[1][2].tag_reg.qe       = reg2hw.tag_258.qe;
  assign rcache_line[1][2].tag_reg.re       = reg2hw.tag_258.re;
  assign rcache_line[1][2].status_reg.status = reg2hw.status_258.q;//status_reg_t'(reg2hw.status_258.q);
  assign rcache_line[1][2].status_reg.qe    = reg2hw.status_258.qe;
  assign rcache_line[1][2].status_reg.re    = reg2hw.status_258.re;


  assign rcache_line[1][3].tag_reg.tag      = reg2hw.tag_259.q;
  assign rcache_line[1][3].tag_reg.qe       = reg2hw.tag_259.qe;
  assign rcache_line[1][3].tag_reg.re       = reg2hw.tag_259.re;
  assign rcache_line[1][3].status_reg.status = reg2hw.status_259.q;//status_reg_t'(reg2hw.status_259.q);
  assign rcache_line[1][3].status_reg.qe    = reg2hw.status_259.qe;
  assign rcache_line[1][3].status_reg.re    = reg2hw.status_259.re;


  assign rcache_line[1][4].tag_reg.tag      = reg2hw.tag_260.q;
  assign rcache_line[1][4].tag_reg.qe       = reg2hw.tag_260.qe;
  assign rcache_line[1][4].tag_reg.re       = reg2hw.tag_260.re;
  assign rcache_line[1][4].status_reg.status = reg2hw.status_260.q;//status_reg_t'(reg2hw.status_260.q);
  assign rcache_line[1][4].status_reg.qe    = reg2hw.status_260.qe;
  assign rcache_line[1][4].status_reg.re    = reg2hw.status_260.re;


  assign rcache_line[1][5].tag_reg.tag      = reg2hw.tag_261.q;
  assign rcache_line[1][5].tag_reg.qe       = reg2hw.tag_261.qe;
  assign rcache_line[1][5].tag_reg.re       = reg2hw.tag_261.re;
  assign rcache_line[1][5].status_reg.status = reg2hw.status_261.q;//status_reg_t'(reg2hw.status_261.q);
  assign rcache_line[1][5].status_reg.qe    = reg2hw.status_261.qe;
  assign rcache_line[1][5].status_reg.re    = reg2hw.status_261.re;


  assign rcache_line[1][6].tag_reg.tag      = reg2hw.tag_262.q;
  assign rcache_line[1][6].tag_reg.qe       = reg2hw.tag_262.qe;
  assign rcache_line[1][6].tag_reg.re       = reg2hw.tag_262.re;
  assign rcache_line[1][6].status_reg.status = reg2hw.status_262.q;//status_reg_t'(reg2hw.status_262.q);
  assign rcache_line[1][6].status_reg.qe    = reg2hw.status_262.qe;
  assign rcache_line[1][6].status_reg.re    = reg2hw.status_262.re;


  assign rcache_line[1][7].tag_reg.tag      = reg2hw.tag_263.q;
  assign rcache_line[1][7].tag_reg.qe       = reg2hw.tag_263.qe;
  assign rcache_line[1][7].tag_reg.re       = reg2hw.tag_263.re;
  assign rcache_line[1][7].status_reg.status = reg2hw.status_263.q;//status_reg_t'(reg2hw.status_263.q);
  assign rcache_line[1][7].status_reg.qe    = reg2hw.status_263.qe;
  assign rcache_line[1][7].status_reg.re    = reg2hw.status_263.re;


  assign rcache_line[1][8].tag_reg.tag      = reg2hw.tag_264.q;
  assign rcache_line[1][8].tag_reg.qe       = reg2hw.tag_264.qe;
  assign rcache_line[1][8].tag_reg.re       = reg2hw.tag_264.re;
  assign rcache_line[1][8].status_reg.status = reg2hw.status_264.q;//status_reg_t'(reg2hw.status_264.q);
  assign rcache_line[1][8].status_reg.qe    = reg2hw.status_264.qe;
  assign rcache_line[1][8].status_reg.re    = reg2hw.status_264.re;


  assign rcache_line[1][9].tag_reg.tag      = reg2hw.tag_265.q;
  assign rcache_line[1][9].tag_reg.qe       = reg2hw.tag_265.qe;
  assign rcache_line[1][9].tag_reg.re       = reg2hw.tag_265.re;
  assign rcache_line[1][9].status_reg.status = reg2hw.status_265.q;//status_reg_t'(reg2hw.status_265.q);
  assign rcache_line[1][9].status_reg.qe    = reg2hw.status_265.qe;
  assign rcache_line[1][9].status_reg.re    = reg2hw.status_265.re;


  assign rcache_line[1][10].tag_reg.tag      = reg2hw.tag_266.q;
  assign rcache_line[1][10].tag_reg.qe       = reg2hw.tag_266.qe;
  assign rcache_line[1][10].tag_reg.re       = reg2hw.tag_266.re;
  assign rcache_line[1][10].status_reg.status = reg2hw.status_266.q;//status_reg_t'(reg2hw.status_266.q);
  assign rcache_line[1][10].status_reg.qe    = reg2hw.status_266.qe;
  assign rcache_line[1][10].status_reg.re    = reg2hw.status_266.re;


  assign rcache_line[1][11].tag_reg.tag      = reg2hw.tag_267.q;
  assign rcache_line[1][11].tag_reg.qe       = reg2hw.tag_267.qe;
  assign rcache_line[1][11].tag_reg.re       = reg2hw.tag_267.re;
  assign rcache_line[1][11].status_reg.status = reg2hw.status_267.q;//status_reg_t'(reg2hw.status_267.q);
  assign rcache_line[1][11].status_reg.qe    = reg2hw.status_267.qe;
  assign rcache_line[1][11].status_reg.re    = reg2hw.status_267.re;


  assign rcache_line[1][12].tag_reg.tag      = reg2hw.tag_268.q;
  assign rcache_line[1][12].tag_reg.qe       = reg2hw.tag_268.qe;
  assign rcache_line[1][12].tag_reg.re       = reg2hw.tag_268.re;
  assign rcache_line[1][12].status_reg.status = reg2hw.status_268.q;//status_reg_t'(reg2hw.status_268.q);
  assign rcache_line[1][12].status_reg.qe    = reg2hw.status_268.qe;
  assign rcache_line[1][12].status_reg.re    = reg2hw.status_268.re;


  assign rcache_line[1][13].tag_reg.tag      = reg2hw.tag_269.q;
  assign rcache_line[1][13].tag_reg.qe       = reg2hw.tag_269.qe;
  assign rcache_line[1][13].tag_reg.re       = reg2hw.tag_269.re;
  assign rcache_line[1][13].status_reg.status = reg2hw.status_269.q;//status_reg_t'(reg2hw.status_269.q);
  assign rcache_line[1][13].status_reg.qe    = reg2hw.status_269.qe;
  assign rcache_line[1][13].status_reg.re    = reg2hw.status_269.re;


  assign rcache_line[1][14].tag_reg.tag      = reg2hw.tag_270.q;
  assign rcache_line[1][14].tag_reg.qe       = reg2hw.tag_270.qe;
  assign rcache_line[1][14].tag_reg.re       = reg2hw.tag_270.re;
  assign rcache_line[1][14].status_reg.status = reg2hw.status_270.q;//status_reg_t'(reg2hw.status_270.q);
  assign rcache_line[1][14].status_reg.qe    = reg2hw.status_270.qe;
  assign rcache_line[1][14].status_reg.re    = reg2hw.status_270.re;


  assign rcache_line[1][15].tag_reg.tag      = reg2hw.tag_271.q;
  assign rcache_line[1][15].tag_reg.qe       = reg2hw.tag_271.qe;
  assign rcache_line[1][15].tag_reg.re       = reg2hw.tag_271.re;
  assign rcache_line[1][15].status_reg.status = reg2hw.status_271.q;//status_reg_t'(reg2hw.status_271.q);
  assign rcache_line[1][15].status_reg.qe    = reg2hw.status_271.qe;
  assign rcache_line[1][15].status_reg.re    = reg2hw.status_271.re;


  assign rcache_line[1][16].tag_reg.tag      = reg2hw.tag_272.q;
  assign rcache_line[1][16].tag_reg.qe       = reg2hw.tag_272.qe;
  assign rcache_line[1][16].tag_reg.re       = reg2hw.tag_272.re;
  assign rcache_line[1][16].status_reg.status = reg2hw.status_272.q;//status_reg_t'(reg2hw.status_272.q);
  assign rcache_line[1][16].status_reg.qe    = reg2hw.status_272.qe;
  assign rcache_line[1][16].status_reg.re    = reg2hw.status_272.re;


  assign rcache_line[1][17].tag_reg.tag      = reg2hw.tag_273.q;
  assign rcache_line[1][17].tag_reg.qe       = reg2hw.tag_273.qe;
  assign rcache_line[1][17].tag_reg.re       = reg2hw.tag_273.re;
  assign rcache_line[1][17].status_reg.status = reg2hw.status_273.q;//status_reg_t'(reg2hw.status_273.q);
  assign rcache_line[1][17].status_reg.qe    = reg2hw.status_273.qe;
  assign rcache_line[1][17].status_reg.re    = reg2hw.status_273.re;


  assign rcache_line[1][18].tag_reg.tag      = reg2hw.tag_274.q;
  assign rcache_line[1][18].tag_reg.qe       = reg2hw.tag_274.qe;
  assign rcache_line[1][18].tag_reg.re       = reg2hw.tag_274.re;
  assign rcache_line[1][18].status_reg.status = reg2hw.status_274.q;//status_reg_t'(reg2hw.status_274.q);
  assign rcache_line[1][18].status_reg.qe    = reg2hw.status_274.qe;
  assign rcache_line[1][18].status_reg.re    = reg2hw.status_274.re;


  assign rcache_line[1][19].tag_reg.tag      = reg2hw.tag_275.q;
  assign rcache_line[1][19].tag_reg.qe       = reg2hw.tag_275.qe;
  assign rcache_line[1][19].tag_reg.re       = reg2hw.tag_275.re;
  assign rcache_line[1][19].status_reg.status = reg2hw.status_275.q;//status_reg_t'(reg2hw.status_275.q);
  assign rcache_line[1][19].status_reg.qe    = reg2hw.status_275.qe;
  assign rcache_line[1][19].status_reg.re    = reg2hw.status_275.re;


  assign rcache_line[1][20].tag_reg.tag      = reg2hw.tag_276.q;
  assign rcache_line[1][20].tag_reg.qe       = reg2hw.tag_276.qe;
  assign rcache_line[1][20].tag_reg.re       = reg2hw.tag_276.re;
  assign rcache_line[1][20].status_reg.status = reg2hw.status_276.q;//status_reg_t'(reg2hw.status_276.q);
  assign rcache_line[1][20].status_reg.qe    = reg2hw.status_276.qe;
  assign rcache_line[1][20].status_reg.re    = reg2hw.status_276.re;


  assign rcache_line[1][21].tag_reg.tag      = reg2hw.tag_277.q;
  assign rcache_line[1][21].tag_reg.qe       = reg2hw.tag_277.qe;
  assign rcache_line[1][21].tag_reg.re       = reg2hw.tag_277.re;
  assign rcache_line[1][21].status_reg.status = reg2hw.status_277.q;//status_reg_t'(reg2hw.status_277.q);
  assign rcache_line[1][21].status_reg.qe    = reg2hw.status_277.qe;
  assign rcache_line[1][21].status_reg.re    = reg2hw.status_277.re;


  assign rcache_line[1][22].tag_reg.tag      = reg2hw.tag_278.q;
  assign rcache_line[1][22].tag_reg.qe       = reg2hw.tag_278.qe;
  assign rcache_line[1][22].tag_reg.re       = reg2hw.tag_278.re;
  assign rcache_line[1][22].status_reg.status = reg2hw.status_278.q;//status_reg_t'(reg2hw.status_278.q);
  assign rcache_line[1][22].status_reg.qe    = reg2hw.status_278.qe;
  assign rcache_line[1][22].status_reg.re    = reg2hw.status_278.re;


  assign rcache_line[1][23].tag_reg.tag      = reg2hw.tag_279.q;
  assign rcache_line[1][23].tag_reg.qe       = reg2hw.tag_279.qe;
  assign rcache_line[1][23].tag_reg.re       = reg2hw.tag_279.re;
  assign rcache_line[1][23].status_reg.status = reg2hw.status_279.q;//status_reg_t'(reg2hw.status_279.q);
  assign rcache_line[1][23].status_reg.qe    = reg2hw.status_279.qe;
  assign rcache_line[1][23].status_reg.re    = reg2hw.status_279.re;


  assign rcache_line[1][24].tag_reg.tag      = reg2hw.tag_280.q;
  assign rcache_line[1][24].tag_reg.qe       = reg2hw.tag_280.qe;
  assign rcache_line[1][24].tag_reg.re       = reg2hw.tag_280.re;
  assign rcache_line[1][24].status_reg.status = reg2hw.status_280.q;//status_reg_t'(reg2hw.status_280.q);
  assign rcache_line[1][24].status_reg.qe    = reg2hw.status_280.qe;
  assign rcache_line[1][24].status_reg.re    = reg2hw.status_280.re;


  assign rcache_line[1][25].tag_reg.tag      = reg2hw.tag_281.q;
  assign rcache_line[1][25].tag_reg.qe       = reg2hw.tag_281.qe;
  assign rcache_line[1][25].tag_reg.re       = reg2hw.tag_281.re;
  assign rcache_line[1][25].status_reg.status = reg2hw.status_281.q;//status_reg_t'(reg2hw.status_281.q);
  assign rcache_line[1][25].status_reg.qe    = reg2hw.status_281.qe;
  assign rcache_line[1][25].status_reg.re    = reg2hw.status_281.re;


  assign rcache_line[1][26].tag_reg.tag      = reg2hw.tag_282.q;
  assign rcache_line[1][26].tag_reg.qe       = reg2hw.tag_282.qe;
  assign rcache_line[1][26].tag_reg.re       = reg2hw.tag_282.re;
  assign rcache_line[1][26].status_reg.status = reg2hw.status_282.q;//status_reg_t'(reg2hw.status_282.q);
  assign rcache_line[1][26].status_reg.qe    = reg2hw.status_282.qe;
  assign rcache_line[1][26].status_reg.re    = reg2hw.status_282.re;


  assign rcache_line[1][27].tag_reg.tag      = reg2hw.tag_283.q;
  assign rcache_line[1][27].tag_reg.qe       = reg2hw.tag_283.qe;
  assign rcache_line[1][27].tag_reg.re       = reg2hw.tag_283.re;
  assign rcache_line[1][27].status_reg.status = reg2hw.status_283.q;//status_reg_t'(reg2hw.status_283.q);
  assign rcache_line[1][27].status_reg.qe    = reg2hw.status_283.qe;
  assign rcache_line[1][27].status_reg.re    = reg2hw.status_283.re;


  assign rcache_line[1][28].tag_reg.tag      = reg2hw.tag_284.q;
  assign rcache_line[1][28].tag_reg.qe       = reg2hw.tag_284.qe;
  assign rcache_line[1][28].tag_reg.re       = reg2hw.tag_284.re;
  assign rcache_line[1][28].status_reg.status = reg2hw.status_284.q;//status_reg_t'(reg2hw.status_284.q);
  assign rcache_line[1][28].status_reg.qe    = reg2hw.status_284.qe;
  assign rcache_line[1][28].status_reg.re    = reg2hw.status_284.re;


  assign rcache_line[1][29].tag_reg.tag      = reg2hw.tag_285.q;
  assign rcache_line[1][29].tag_reg.qe       = reg2hw.tag_285.qe;
  assign rcache_line[1][29].tag_reg.re       = reg2hw.tag_285.re;
  assign rcache_line[1][29].status_reg.status = reg2hw.status_285.q;//status_reg_t'(reg2hw.status_285.q);
  assign rcache_line[1][29].status_reg.qe    = reg2hw.status_285.qe;
  assign rcache_line[1][29].status_reg.re    = reg2hw.status_285.re;


  assign rcache_line[1][30].tag_reg.tag      = reg2hw.tag_286.q;
  assign rcache_line[1][30].tag_reg.qe       = reg2hw.tag_286.qe;
  assign rcache_line[1][30].tag_reg.re       = reg2hw.tag_286.re;
  assign rcache_line[1][30].status_reg.status = reg2hw.status_286.q;//status_reg_t'(reg2hw.status_286.q);
  assign rcache_line[1][30].status_reg.qe    = reg2hw.status_286.qe;
  assign rcache_line[1][30].status_reg.re    = reg2hw.status_286.re;


  assign rcache_line[1][31].tag_reg.tag      = reg2hw.tag_287.q;
  assign rcache_line[1][31].tag_reg.qe       = reg2hw.tag_287.qe;
  assign rcache_line[1][31].tag_reg.re       = reg2hw.tag_287.re;
  assign rcache_line[1][31].status_reg.status = reg2hw.status_287.q;//status_reg_t'(reg2hw.status_287.q);
  assign rcache_line[1][31].status_reg.qe    = reg2hw.status_287.qe;
  assign rcache_line[1][31].status_reg.re    = reg2hw.status_287.re;


  assign rcache_line[1][32].tag_reg.tag      = reg2hw.tag_288.q;
  assign rcache_line[1][32].tag_reg.qe       = reg2hw.tag_288.qe;
  assign rcache_line[1][32].tag_reg.re       = reg2hw.tag_288.re;
  assign rcache_line[1][32].status_reg.status = reg2hw.status_288.q;//status_reg_t'(reg2hw.status_288.q);
  assign rcache_line[1][32].status_reg.qe    = reg2hw.status_288.qe;
  assign rcache_line[1][32].status_reg.re    = reg2hw.status_288.re;


  assign rcache_line[1][33].tag_reg.tag      = reg2hw.tag_289.q;
  assign rcache_line[1][33].tag_reg.qe       = reg2hw.tag_289.qe;
  assign rcache_line[1][33].tag_reg.re       = reg2hw.tag_289.re;
  assign rcache_line[1][33].status_reg.status = reg2hw.status_289.q;//status_reg_t'(reg2hw.status_289.q);
  assign rcache_line[1][33].status_reg.qe    = reg2hw.status_289.qe;
  assign rcache_line[1][33].status_reg.re    = reg2hw.status_289.re;


  assign rcache_line[1][34].tag_reg.tag      = reg2hw.tag_290.q;
  assign rcache_line[1][34].tag_reg.qe       = reg2hw.tag_290.qe;
  assign rcache_line[1][34].tag_reg.re       = reg2hw.tag_290.re;
  assign rcache_line[1][34].status_reg.status = reg2hw.status_290.q;//status_reg_t'(reg2hw.status_290.q);
  assign rcache_line[1][34].status_reg.qe    = reg2hw.status_290.qe;
  assign rcache_line[1][34].status_reg.re    = reg2hw.status_290.re;


  assign rcache_line[1][35].tag_reg.tag      = reg2hw.tag_291.q;
  assign rcache_line[1][35].tag_reg.qe       = reg2hw.tag_291.qe;
  assign rcache_line[1][35].tag_reg.re       = reg2hw.tag_291.re;
  assign rcache_line[1][35].status_reg.status = reg2hw.status_291.q;//status_reg_t'(reg2hw.status_291.q);
  assign rcache_line[1][35].status_reg.qe    = reg2hw.status_291.qe;
  assign rcache_line[1][35].status_reg.re    = reg2hw.status_291.re;


  assign rcache_line[1][36].tag_reg.tag      = reg2hw.tag_292.q;
  assign rcache_line[1][36].tag_reg.qe       = reg2hw.tag_292.qe;
  assign rcache_line[1][36].tag_reg.re       = reg2hw.tag_292.re;
  assign rcache_line[1][36].status_reg.status = reg2hw.status_292.q;//status_reg_t'(reg2hw.status_292.q);
  assign rcache_line[1][36].status_reg.qe    = reg2hw.status_292.qe;
  assign rcache_line[1][36].status_reg.re    = reg2hw.status_292.re;


  assign rcache_line[1][37].tag_reg.tag      = reg2hw.tag_293.q;
  assign rcache_line[1][37].tag_reg.qe       = reg2hw.tag_293.qe;
  assign rcache_line[1][37].tag_reg.re       = reg2hw.tag_293.re;
  assign rcache_line[1][37].status_reg.status = reg2hw.status_293.q;//status_reg_t'(reg2hw.status_293.q);
  assign rcache_line[1][37].status_reg.qe    = reg2hw.status_293.qe;
  assign rcache_line[1][37].status_reg.re    = reg2hw.status_293.re;


  assign rcache_line[1][38].tag_reg.tag      = reg2hw.tag_294.q;
  assign rcache_line[1][38].tag_reg.qe       = reg2hw.tag_294.qe;
  assign rcache_line[1][38].tag_reg.re       = reg2hw.tag_294.re;
  assign rcache_line[1][38].status_reg.status = reg2hw.status_294.q;//status_reg_t'(reg2hw.status_294.q);
  assign rcache_line[1][38].status_reg.qe    = reg2hw.status_294.qe;
  assign rcache_line[1][38].status_reg.re    = reg2hw.status_294.re;


  assign rcache_line[1][39].tag_reg.tag      = reg2hw.tag_295.q;
  assign rcache_line[1][39].tag_reg.qe       = reg2hw.tag_295.qe;
  assign rcache_line[1][39].tag_reg.re       = reg2hw.tag_295.re;
  assign rcache_line[1][39].status_reg.status = reg2hw.status_295.q;//status_reg_t'(reg2hw.status_295.q);
  assign rcache_line[1][39].status_reg.qe    = reg2hw.status_295.qe;
  assign rcache_line[1][39].status_reg.re    = reg2hw.status_295.re;


  assign rcache_line[1][40].tag_reg.tag      = reg2hw.tag_296.q;
  assign rcache_line[1][40].tag_reg.qe       = reg2hw.tag_296.qe;
  assign rcache_line[1][40].tag_reg.re       = reg2hw.tag_296.re;
  assign rcache_line[1][40].status_reg.status = reg2hw.status_296.q;//status_reg_t'(reg2hw.status_296.q);
  assign rcache_line[1][40].status_reg.qe    = reg2hw.status_296.qe;
  assign rcache_line[1][40].status_reg.re    = reg2hw.status_296.re;


  assign rcache_line[1][41].tag_reg.tag      = reg2hw.tag_297.q;
  assign rcache_line[1][41].tag_reg.qe       = reg2hw.tag_297.qe;
  assign rcache_line[1][41].tag_reg.re       = reg2hw.tag_297.re;
  assign rcache_line[1][41].status_reg.status = reg2hw.status_297.q;//status_reg_t'(reg2hw.status_297.q);
  assign rcache_line[1][41].status_reg.qe    = reg2hw.status_297.qe;
  assign rcache_line[1][41].status_reg.re    = reg2hw.status_297.re;


  assign rcache_line[1][42].tag_reg.tag      = reg2hw.tag_298.q;
  assign rcache_line[1][42].tag_reg.qe       = reg2hw.tag_298.qe;
  assign rcache_line[1][42].tag_reg.re       = reg2hw.tag_298.re;
  assign rcache_line[1][42].status_reg.status = reg2hw.status_298.q;//status_reg_t'(reg2hw.status_298.q);
  assign rcache_line[1][42].status_reg.qe    = reg2hw.status_298.qe;
  assign rcache_line[1][42].status_reg.re    = reg2hw.status_298.re;


  assign rcache_line[1][43].tag_reg.tag      = reg2hw.tag_299.q;
  assign rcache_line[1][43].tag_reg.qe       = reg2hw.tag_299.qe;
  assign rcache_line[1][43].tag_reg.re       = reg2hw.tag_299.re;
  assign rcache_line[1][43].status_reg.status = reg2hw.status_299.q;//status_reg_t'(reg2hw.status_299.q);
  assign rcache_line[1][43].status_reg.qe    = reg2hw.status_299.qe;
  assign rcache_line[1][43].status_reg.re    = reg2hw.status_299.re;


  assign rcache_line[1][44].tag_reg.tag      = reg2hw.tag_300.q;
  assign rcache_line[1][44].tag_reg.qe       = reg2hw.tag_300.qe;
  assign rcache_line[1][44].tag_reg.re       = reg2hw.tag_300.re;
  assign rcache_line[1][44].status_reg.status = reg2hw.status_300.q;//status_reg_t'(reg2hw.status_300.q);
  assign rcache_line[1][44].status_reg.qe    = reg2hw.status_300.qe;
  assign rcache_line[1][44].status_reg.re    = reg2hw.status_300.re;


  assign rcache_line[1][45].tag_reg.tag      = reg2hw.tag_301.q;
  assign rcache_line[1][45].tag_reg.qe       = reg2hw.tag_301.qe;
  assign rcache_line[1][45].tag_reg.re       = reg2hw.tag_301.re;
  assign rcache_line[1][45].status_reg.status = reg2hw.status_301.q;//status_reg_t'(reg2hw.status_301.q);
  assign rcache_line[1][45].status_reg.qe    = reg2hw.status_301.qe;
  assign rcache_line[1][45].status_reg.re    = reg2hw.status_301.re;


  assign rcache_line[1][46].tag_reg.tag      = reg2hw.tag_302.q;
  assign rcache_line[1][46].tag_reg.qe       = reg2hw.tag_302.qe;
  assign rcache_line[1][46].tag_reg.re       = reg2hw.tag_302.re;
  assign rcache_line[1][46].status_reg.status = reg2hw.status_302.q;//status_reg_t'(reg2hw.status_302.q);
  assign rcache_line[1][46].status_reg.qe    = reg2hw.status_302.qe;
  assign rcache_line[1][46].status_reg.re    = reg2hw.status_302.re;


  assign rcache_line[1][47].tag_reg.tag      = reg2hw.tag_303.q;
  assign rcache_line[1][47].tag_reg.qe       = reg2hw.tag_303.qe;
  assign rcache_line[1][47].tag_reg.re       = reg2hw.tag_303.re;
  assign rcache_line[1][47].status_reg.status = reg2hw.status_303.q;//status_reg_t'(reg2hw.status_303.q);
  assign rcache_line[1][47].status_reg.qe    = reg2hw.status_303.qe;
  assign rcache_line[1][47].status_reg.re    = reg2hw.status_303.re;


  assign rcache_line[1][48].tag_reg.tag      = reg2hw.tag_304.q;
  assign rcache_line[1][48].tag_reg.qe       = reg2hw.tag_304.qe;
  assign rcache_line[1][48].tag_reg.re       = reg2hw.tag_304.re;
  assign rcache_line[1][48].status_reg.status = reg2hw.status_304.q;//status_reg_t'(reg2hw.status_304.q);
  assign rcache_line[1][48].status_reg.qe    = reg2hw.status_304.qe;
  assign rcache_line[1][48].status_reg.re    = reg2hw.status_304.re;


  assign rcache_line[1][49].tag_reg.tag      = reg2hw.tag_305.q;
  assign rcache_line[1][49].tag_reg.qe       = reg2hw.tag_305.qe;
  assign rcache_line[1][49].tag_reg.re       = reg2hw.tag_305.re;
  assign rcache_line[1][49].status_reg.status = reg2hw.status_305.q;//status_reg_t'(reg2hw.status_305.q);
  assign rcache_line[1][49].status_reg.qe    = reg2hw.status_305.qe;
  assign rcache_line[1][49].status_reg.re    = reg2hw.status_305.re;


  assign rcache_line[1][50].tag_reg.tag      = reg2hw.tag_306.q;
  assign rcache_line[1][50].tag_reg.qe       = reg2hw.tag_306.qe;
  assign rcache_line[1][50].tag_reg.re       = reg2hw.tag_306.re;
  assign rcache_line[1][50].status_reg.status = reg2hw.status_306.q;//status_reg_t'(reg2hw.status_306.q);
  assign rcache_line[1][50].status_reg.qe    = reg2hw.status_306.qe;
  assign rcache_line[1][50].status_reg.re    = reg2hw.status_306.re;


  assign rcache_line[1][51].tag_reg.tag      = reg2hw.tag_307.q;
  assign rcache_line[1][51].tag_reg.qe       = reg2hw.tag_307.qe;
  assign rcache_line[1][51].tag_reg.re       = reg2hw.tag_307.re;
  assign rcache_line[1][51].status_reg.status = reg2hw.status_307.q;//status_reg_t'(reg2hw.status_307.q);
  assign rcache_line[1][51].status_reg.qe    = reg2hw.status_307.qe;
  assign rcache_line[1][51].status_reg.re    = reg2hw.status_307.re;


  assign rcache_line[1][52].tag_reg.tag      = reg2hw.tag_308.q;
  assign rcache_line[1][52].tag_reg.qe       = reg2hw.tag_308.qe;
  assign rcache_line[1][52].tag_reg.re       = reg2hw.tag_308.re;
  assign rcache_line[1][52].status_reg.status = reg2hw.status_308.q;//status_reg_t'(reg2hw.status_308.q);
  assign rcache_line[1][52].status_reg.qe    = reg2hw.status_308.qe;
  assign rcache_line[1][52].status_reg.re    = reg2hw.status_308.re;


  assign rcache_line[1][53].tag_reg.tag      = reg2hw.tag_309.q;
  assign rcache_line[1][53].tag_reg.qe       = reg2hw.tag_309.qe;
  assign rcache_line[1][53].tag_reg.re       = reg2hw.tag_309.re;
  assign rcache_line[1][53].status_reg.status = reg2hw.status_309.q;//status_reg_t'(reg2hw.status_309.q);
  assign rcache_line[1][53].status_reg.qe    = reg2hw.status_309.qe;
  assign rcache_line[1][53].status_reg.re    = reg2hw.status_309.re;


  assign rcache_line[1][54].tag_reg.tag      = reg2hw.tag_310.q;
  assign rcache_line[1][54].tag_reg.qe       = reg2hw.tag_310.qe;
  assign rcache_line[1][54].tag_reg.re       = reg2hw.tag_310.re;
  assign rcache_line[1][54].status_reg.status = reg2hw.status_310.q;//status_reg_t'(reg2hw.status_310.q);
  assign rcache_line[1][54].status_reg.qe    = reg2hw.status_310.qe;
  assign rcache_line[1][54].status_reg.re    = reg2hw.status_310.re;


  assign rcache_line[1][55].tag_reg.tag      = reg2hw.tag_311.q;
  assign rcache_line[1][55].tag_reg.qe       = reg2hw.tag_311.qe;
  assign rcache_line[1][55].tag_reg.re       = reg2hw.tag_311.re;
  assign rcache_line[1][55].status_reg.status = reg2hw.status_311.q;//status_reg_t'(reg2hw.status_311.q);
  assign rcache_line[1][55].status_reg.qe    = reg2hw.status_311.qe;
  assign rcache_line[1][55].status_reg.re    = reg2hw.status_311.re;


  assign rcache_line[1][56].tag_reg.tag      = reg2hw.tag_312.q;
  assign rcache_line[1][56].tag_reg.qe       = reg2hw.tag_312.qe;
  assign rcache_line[1][56].tag_reg.re       = reg2hw.tag_312.re;
  assign rcache_line[1][56].status_reg.status = reg2hw.status_312.q;//status_reg_t'(reg2hw.status_312.q);
  assign rcache_line[1][56].status_reg.qe    = reg2hw.status_312.qe;
  assign rcache_line[1][56].status_reg.re    = reg2hw.status_312.re;


  assign rcache_line[1][57].tag_reg.tag      = reg2hw.tag_313.q;
  assign rcache_line[1][57].tag_reg.qe       = reg2hw.tag_313.qe;
  assign rcache_line[1][57].tag_reg.re       = reg2hw.tag_313.re;
  assign rcache_line[1][57].status_reg.status = reg2hw.status_313.q;//status_reg_t'(reg2hw.status_313.q);
  assign rcache_line[1][57].status_reg.qe    = reg2hw.status_313.qe;
  assign rcache_line[1][57].status_reg.re    = reg2hw.status_313.re;


  assign rcache_line[1][58].tag_reg.tag      = reg2hw.tag_314.q;
  assign rcache_line[1][58].tag_reg.qe       = reg2hw.tag_314.qe;
  assign rcache_line[1][58].tag_reg.re       = reg2hw.tag_314.re;
  assign rcache_line[1][58].status_reg.status = reg2hw.status_314.q;//status_reg_t'(reg2hw.status_314.q);
  assign rcache_line[1][58].status_reg.qe    = reg2hw.status_314.qe;
  assign rcache_line[1][58].status_reg.re    = reg2hw.status_314.re;


  assign rcache_line[1][59].tag_reg.tag      = reg2hw.tag_315.q;
  assign rcache_line[1][59].tag_reg.qe       = reg2hw.tag_315.qe;
  assign rcache_line[1][59].tag_reg.re       = reg2hw.tag_315.re;
  assign rcache_line[1][59].status_reg.status = reg2hw.status_315.q;//status_reg_t'(reg2hw.status_315.q);
  assign rcache_line[1][59].status_reg.qe    = reg2hw.status_315.qe;
  assign rcache_line[1][59].status_reg.re    = reg2hw.status_315.re;


  assign rcache_line[1][60].tag_reg.tag      = reg2hw.tag_316.q;
  assign rcache_line[1][60].tag_reg.qe       = reg2hw.tag_316.qe;
  assign rcache_line[1][60].tag_reg.re       = reg2hw.tag_316.re;
  assign rcache_line[1][60].status_reg.status = reg2hw.status_316.q;//status_reg_t'(reg2hw.status_316.q);
  assign rcache_line[1][60].status_reg.qe    = reg2hw.status_316.qe;
  assign rcache_line[1][60].status_reg.re    = reg2hw.status_316.re;


  assign rcache_line[1][61].tag_reg.tag      = reg2hw.tag_317.q;
  assign rcache_line[1][61].tag_reg.qe       = reg2hw.tag_317.qe;
  assign rcache_line[1][61].tag_reg.re       = reg2hw.tag_317.re;
  assign rcache_line[1][61].status_reg.status = reg2hw.status_317.q;//status_reg_t'(reg2hw.status_317.q);
  assign rcache_line[1][61].status_reg.qe    = reg2hw.status_317.qe;
  assign rcache_line[1][61].status_reg.re    = reg2hw.status_317.re;


  assign rcache_line[1][62].tag_reg.tag      = reg2hw.tag_318.q;
  assign rcache_line[1][62].tag_reg.qe       = reg2hw.tag_318.qe;
  assign rcache_line[1][62].tag_reg.re       = reg2hw.tag_318.re;
  assign rcache_line[1][62].status_reg.status = reg2hw.status_318.q;//status_reg_t'(reg2hw.status_318.q);
  assign rcache_line[1][62].status_reg.qe    = reg2hw.status_318.qe;
  assign rcache_line[1][62].status_reg.re    = reg2hw.status_318.re;


  assign rcache_line[1][63].tag_reg.tag      = reg2hw.tag_319.q;
  assign rcache_line[1][63].tag_reg.qe       = reg2hw.tag_319.qe;
  assign rcache_line[1][63].tag_reg.re       = reg2hw.tag_319.re;
  assign rcache_line[1][63].status_reg.status = reg2hw.status_319.q;//status_reg_t'(reg2hw.status_319.q);
  assign rcache_line[1][63].status_reg.qe    = reg2hw.status_319.qe;
  assign rcache_line[1][63].status_reg.re    = reg2hw.status_319.re;


  assign rcache_line[1][64].tag_reg.tag      = reg2hw.tag_320.q;
  assign rcache_line[1][64].tag_reg.qe       = reg2hw.tag_320.qe;
  assign rcache_line[1][64].tag_reg.re       = reg2hw.tag_320.re;
  assign rcache_line[1][64].status_reg.status = reg2hw.status_320.q;//status_reg_t'(reg2hw.status_320.q);
  assign rcache_line[1][64].status_reg.qe    = reg2hw.status_320.qe;
  assign rcache_line[1][64].status_reg.re    = reg2hw.status_320.re;


  assign rcache_line[1][65].tag_reg.tag      = reg2hw.tag_321.q;
  assign rcache_line[1][65].tag_reg.qe       = reg2hw.tag_321.qe;
  assign rcache_line[1][65].tag_reg.re       = reg2hw.tag_321.re;
  assign rcache_line[1][65].status_reg.status = reg2hw.status_321.q;//status_reg_t'(reg2hw.status_321.q);
  assign rcache_line[1][65].status_reg.qe    = reg2hw.status_321.qe;
  assign rcache_line[1][65].status_reg.re    = reg2hw.status_321.re;


  assign rcache_line[1][66].tag_reg.tag      = reg2hw.tag_322.q;
  assign rcache_line[1][66].tag_reg.qe       = reg2hw.tag_322.qe;
  assign rcache_line[1][66].tag_reg.re       = reg2hw.tag_322.re;
  assign rcache_line[1][66].status_reg.status = reg2hw.status_322.q;//status_reg_t'(reg2hw.status_322.q);
  assign rcache_line[1][66].status_reg.qe    = reg2hw.status_322.qe;
  assign rcache_line[1][66].status_reg.re    = reg2hw.status_322.re;


  assign rcache_line[1][67].tag_reg.tag      = reg2hw.tag_323.q;
  assign rcache_line[1][67].tag_reg.qe       = reg2hw.tag_323.qe;
  assign rcache_line[1][67].tag_reg.re       = reg2hw.tag_323.re;
  assign rcache_line[1][67].status_reg.status = reg2hw.status_323.q;//status_reg_t'(reg2hw.status_323.q);
  assign rcache_line[1][67].status_reg.qe    = reg2hw.status_323.qe;
  assign rcache_line[1][67].status_reg.re    = reg2hw.status_323.re;


  assign rcache_line[1][68].tag_reg.tag      = reg2hw.tag_324.q;
  assign rcache_line[1][68].tag_reg.qe       = reg2hw.tag_324.qe;
  assign rcache_line[1][68].tag_reg.re       = reg2hw.tag_324.re;
  assign rcache_line[1][68].status_reg.status = reg2hw.status_324.q;//status_reg_t'(reg2hw.status_324.q);
  assign rcache_line[1][68].status_reg.qe    = reg2hw.status_324.qe;
  assign rcache_line[1][68].status_reg.re    = reg2hw.status_324.re;


  assign rcache_line[1][69].tag_reg.tag      = reg2hw.tag_325.q;
  assign rcache_line[1][69].tag_reg.qe       = reg2hw.tag_325.qe;
  assign rcache_line[1][69].tag_reg.re       = reg2hw.tag_325.re;
  assign rcache_line[1][69].status_reg.status = reg2hw.status_325.q;//status_reg_t'(reg2hw.status_325.q);
  assign rcache_line[1][69].status_reg.qe    = reg2hw.status_325.qe;
  assign rcache_line[1][69].status_reg.re    = reg2hw.status_325.re;


  assign rcache_line[1][70].tag_reg.tag      = reg2hw.tag_326.q;
  assign rcache_line[1][70].tag_reg.qe       = reg2hw.tag_326.qe;
  assign rcache_line[1][70].tag_reg.re       = reg2hw.tag_326.re;
  assign rcache_line[1][70].status_reg.status = reg2hw.status_326.q;//status_reg_t'(reg2hw.status_326.q);
  assign rcache_line[1][70].status_reg.qe    = reg2hw.status_326.qe;
  assign rcache_line[1][70].status_reg.re    = reg2hw.status_326.re;


  assign rcache_line[1][71].tag_reg.tag      = reg2hw.tag_327.q;
  assign rcache_line[1][71].tag_reg.qe       = reg2hw.tag_327.qe;
  assign rcache_line[1][71].tag_reg.re       = reg2hw.tag_327.re;
  assign rcache_line[1][71].status_reg.status = reg2hw.status_327.q;//status_reg_t'(reg2hw.status_327.q);
  assign rcache_line[1][71].status_reg.qe    = reg2hw.status_327.qe;
  assign rcache_line[1][71].status_reg.re    = reg2hw.status_327.re;


  assign rcache_line[1][72].tag_reg.tag      = reg2hw.tag_328.q;
  assign rcache_line[1][72].tag_reg.qe       = reg2hw.tag_328.qe;
  assign rcache_line[1][72].tag_reg.re       = reg2hw.tag_328.re;
  assign rcache_line[1][72].status_reg.status = reg2hw.status_328.q;//status_reg_t'(reg2hw.status_328.q);
  assign rcache_line[1][72].status_reg.qe    = reg2hw.status_328.qe;
  assign rcache_line[1][72].status_reg.re    = reg2hw.status_328.re;


  assign rcache_line[1][73].tag_reg.tag      = reg2hw.tag_329.q;
  assign rcache_line[1][73].tag_reg.qe       = reg2hw.tag_329.qe;
  assign rcache_line[1][73].tag_reg.re       = reg2hw.tag_329.re;
  assign rcache_line[1][73].status_reg.status = reg2hw.status_329.q;//status_reg_t'(reg2hw.status_329.q);
  assign rcache_line[1][73].status_reg.qe    = reg2hw.status_329.qe;
  assign rcache_line[1][73].status_reg.re    = reg2hw.status_329.re;


  assign rcache_line[1][74].tag_reg.tag      = reg2hw.tag_330.q;
  assign rcache_line[1][74].tag_reg.qe       = reg2hw.tag_330.qe;
  assign rcache_line[1][74].tag_reg.re       = reg2hw.tag_330.re;
  assign rcache_line[1][74].status_reg.status = reg2hw.status_330.q;//status_reg_t'(reg2hw.status_330.q);
  assign rcache_line[1][74].status_reg.qe    = reg2hw.status_330.qe;
  assign rcache_line[1][74].status_reg.re    = reg2hw.status_330.re;


  assign rcache_line[1][75].tag_reg.tag      = reg2hw.tag_331.q;
  assign rcache_line[1][75].tag_reg.qe       = reg2hw.tag_331.qe;
  assign rcache_line[1][75].tag_reg.re       = reg2hw.tag_331.re;
  assign rcache_line[1][75].status_reg.status = reg2hw.status_331.q;//status_reg_t'(reg2hw.status_331.q);
  assign rcache_line[1][75].status_reg.qe    = reg2hw.status_331.qe;
  assign rcache_line[1][75].status_reg.re    = reg2hw.status_331.re;


  assign rcache_line[1][76].tag_reg.tag      = reg2hw.tag_332.q;
  assign rcache_line[1][76].tag_reg.qe       = reg2hw.tag_332.qe;
  assign rcache_line[1][76].tag_reg.re       = reg2hw.tag_332.re;
  assign rcache_line[1][76].status_reg.status = reg2hw.status_332.q;//status_reg_t'(reg2hw.status_332.q);
  assign rcache_line[1][76].status_reg.qe    = reg2hw.status_332.qe;
  assign rcache_line[1][76].status_reg.re    = reg2hw.status_332.re;


  assign rcache_line[1][77].tag_reg.tag      = reg2hw.tag_333.q;
  assign rcache_line[1][77].tag_reg.qe       = reg2hw.tag_333.qe;
  assign rcache_line[1][77].tag_reg.re       = reg2hw.tag_333.re;
  assign rcache_line[1][77].status_reg.status = reg2hw.status_333.q;//status_reg_t'(reg2hw.status_333.q);
  assign rcache_line[1][77].status_reg.qe    = reg2hw.status_333.qe;
  assign rcache_line[1][77].status_reg.re    = reg2hw.status_333.re;


  assign rcache_line[1][78].tag_reg.tag      = reg2hw.tag_334.q;
  assign rcache_line[1][78].tag_reg.qe       = reg2hw.tag_334.qe;
  assign rcache_line[1][78].tag_reg.re       = reg2hw.tag_334.re;
  assign rcache_line[1][78].status_reg.status = reg2hw.status_334.q;//status_reg_t'(reg2hw.status_334.q);
  assign rcache_line[1][78].status_reg.qe    = reg2hw.status_334.qe;
  assign rcache_line[1][78].status_reg.re    = reg2hw.status_334.re;


  assign rcache_line[1][79].tag_reg.tag      = reg2hw.tag_335.q;
  assign rcache_line[1][79].tag_reg.qe       = reg2hw.tag_335.qe;
  assign rcache_line[1][79].tag_reg.re       = reg2hw.tag_335.re;
  assign rcache_line[1][79].status_reg.status = reg2hw.status_335.q;//status_reg_t'(reg2hw.status_335.q);
  assign rcache_line[1][79].status_reg.qe    = reg2hw.status_335.qe;
  assign rcache_line[1][79].status_reg.re    = reg2hw.status_335.re;


  assign rcache_line[1][80].tag_reg.tag      = reg2hw.tag_336.q;
  assign rcache_line[1][80].tag_reg.qe       = reg2hw.tag_336.qe;
  assign rcache_line[1][80].tag_reg.re       = reg2hw.tag_336.re;
  assign rcache_line[1][80].status_reg.status = reg2hw.status_336.q;//status_reg_t'(reg2hw.status_336.q);
  assign rcache_line[1][80].status_reg.qe    = reg2hw.status_336.qe;
  assign rcache_line[1][80].status_reg.re    = reg2hw.status_336.re;


  assign rcache_line[1][81].tag_reg.tag      = reg2hw.tag_337.q;
  assign rcache_line[1][81].tag_reg.qe       = reg2hw.tag_337.qe;
  assign rcache_line[1][81].tag_reg.re       = reg2hw.tag_337.re;
  assign rcache_line[1][81].status_reg.status = reg2hw.status_337.q;//status_reg_t'(reg2hw.status_337.q);
  assign rcache_line[1][81].status_reg.qe    = reg2hw.status_337.qe;
  assign rcache_line[1][81].status_reg.re    = reg2hw.status_337.re;


  assign rcache_line[1][82].tag_reg.tag      = reg2hw.tag_338.q;
  assign rcache_line[1][82].tag_reg.qe       = reg2hw.tag_338.qe;
  assign rcache_line[1][82].tag_reg.re       = reg2hw.tag_338.re;
  assign rcache_line[1][82].status_reg.status = reg2hw.status_338.q;//status_reg_t'(reg2hw.status_338.q);
  assign rcache_line[1][82].status_reg.qe    = reg2hw.status_338.qe;
  assign rcache_line[1][82].status_reg.re    = reg2hw.status_338.re;


  assign rcache_line[1][83].tag_reg.tag      = reg2hw.tag_339.q;
  assign rcache_line[1][83].tag_reg.qe       = reg2hw.tag_339.qe;
  assign rcache_line[1][83].tag_reg.re       = reg2hw.tag_339.re;
  assign rcache_line[1][83].status_reg.status = reg2hw.status_339.q;//status_reg_t'(reg2hw.status_339.q);
  assign rcache_line[1][83].status_reg.qe    = reg2hw.status_339.qe;
  assign rcache_line[1][83].status_reg.re    = reg2hw.status_339.re;


  assign rcache_line[1][84].tag_reg.tag      = reg2hw.tag_340.q;
  assign rcache_line[1][84].tag_reg.qe       = reg2hw.tag_340.qe;
  assign rcache_line[1][84].tag_reg.re       = reg2hw.tag_340.re;
  assign rcache_line[1][84].status_reg.status = reg2hw.status_340.q;//status_reg_t'(reg2hw.status_340.q);
  assign rcache_line[1][84].status_reg.qe    = reg2hw.status_340.qe;
  assign rcache_line[1][84].status_reg.re    = reg2hw.status_340.re;


  assign rcache_line[1][85].tag_reg.tag      = reg2hw.tag_341.q;
  assign rcache_line[1][85].tag_reg.qe       = reg2hw.tag_341.qe;
  assign rcache_line[1][85].tag_reg.re       = reg2hw.tag_341.re;
  assign rcache_line[1][85].status_reg.status = reg2hw.status_341.q;//status_reg_t'(reg2hw.status_341.q);
  assign rcache_line[1][85].status_reg.qe    = reg2hw.status_341.qe;
  assign rcache_line[1][85].status_reg.re    = reg2hw.status_341.re;


  assign rcache_line[1][86].tag_reg.tag      = reg2hw.tag_342.q;
  assign rcache_line[1][86].tag_reg.qe       = reg2hw.tag_342.qe;
  assign rcache_line[1][86].tag_reg.re       = reg2hw.tag_342.re;
  assign rcache_line[1][86].status_reg.status = reg2hw.status_342.q;//status_reg_t'(reg2hw.status_342.q);
  assign rcache_line[1][86].status_reg.qe    = reg2hw.status_342.qe;
  assign rcache_line[1][86].status_reg.re    = reg2hw.status_342.re;


  assign rcache_line[1][87].tag_reg.tag      = reg2hw.tag_343.q;
  assign rcache_line[1][87].tag_reg.qe       = reg2hw.tag_343.qe;
  assign rcache_line[1][87].tag_reg.re       = reg2hw.tag_343.re;
  assign rcache_line[1][87].status_reg.status = reg2hw.status_343.q;//status_reg_t'(reg2hw.status_343.q);
  assign rcache_line[1][87].status_reg.qe    = reg2hw.status_343.qe;
  assign rcache_line[1][87].status_reg.re    = reg2hw.status_343.re;


  assign rcache_line[1][88].tag_reg.tag      = reg2hw.tag_344.q;
  assign rcache_line[1][88].tag_reg.qe       = reg2hw.tag_344.qe;
  assign rcache_line[1][88].tag_reg.re       = reg2hw.tag_344.re;
  assign rcache_line[1][88].status_reg.status = reg2hw.status_344.q;//status_reg_t'(reg2hw.status_344.q);
  assign rcache_line[1][88].status_reg.qe    = reg2hw.status_344.qe;
  assign rcache_line[1][88].status_reg.re    = reg2hw.status_344.re;


  assign rcache_line[1][89].tag_reg.tag      = reg2hw.tag_345.q;
  assign rcache_line[1][89].tag_reg.qe       = reg2hw.tag_345.qe;
  assign rcache_line[1][89].tag_reg.re       = reg2hw.tag_345.re;
  assign rcache_line[1][89].status_reg.status = reg2hw.status_345.q;//status_reg_t'(reg2hw.status_345.q);
  assign rcache_line[1][89].status_reg.qe    = reg2hw.status_345.qe;
  assign rcache_line[1][89].status_reg.re    = reg2hw.status_345.re;


  assign rcache_line[1][90].tag_reg.tag      = reg2hw.tag_346.q;
  assign rcache_line[1][90].tag_reg.qe       = reg2hw.tag_346.qe;
  assign rcache_line[1][90].tag_reg.re       = reg2hw.tag_346.re;
  assign rcache_line[1][90].status_reg.status = reg2hw.status_346.q;//status_reg_t'(reg2hw.status_346.q);
  assign rcache_line[1][90].status_reg.qe    = reg2hw.status_346.qe;
  assign rcache_line[1][90].status_reg.re    = reg2hw.status_346.re;


  assign rcache_line[1][91].tag_reg.tag      = reg2hw.tag_347.q;
  assign rcache_line[1][91].tag_reg.qe       = reg2hw.tag_347.qe;
  assign rcache_line[1][91].tag_reg.re       = reg2hw.tag_347.re;
  assign rcache_line[1][91].status_reg.status = reg2hw.status_347.q;//status_reg_t'(reg2hw.status_347.q);
  assign rcache_line[1][91].status_reg.qe    = reg2hw.status_347.qe;
  assign rcache_line[1][91].status_reg.re    = reg2hw.status_347.re;


  assign rcache_line[1][92].tag_reg.tag      = reg2hw.tag_348.q;
  assign rcache_line[1][92].tag_reg.qe       = reg2hw.tag_348.qe;
  assign rcache_line[1][92].tag_reg.re       = reg2hw.tag_348.re;
  assign rcache_line[1][92].status_reg.status = reg2hw.status_348.q;//status_reg_t'(reg2hw.status_348.q);
  assign rcache_line[1][92].status_reg.qe    = reg2hw.status_348.qe;
  assign rcache_line[1][92].status_reg.re    = reg2hw.status_348.re;


  assign rcache_line[1][93].tag_reg.tag      = reg2hw.tag_349.q;
  assign rcache_line[1][93].tag_reg.qe       = reg2hw.tag_349.qe;
  assign rcache_line[1][93].tag_reg.re       = reg2hw.tag_349.re;
  assign rcache_line[1][93].status_reg.status = reg2hw.status_349.q;//status_reg_t'(reg2hw.status_349.q);
  assign rcache_line[1][93].status_reg.qe    = reg2hw.status_349.qe;
  assign rcache_line[1][93].status_reg.re    = reg2hw.status_349.re;


  assign rcache_line[1][94].tag_reg.tag      = reg2hw.tag_350.q;
  assign rcache_line[1][94].tag_reg.qe       = reg2hw.tag_350.qe;
  assign rcache_line[1][94].tag_reg.re       = reg2hw.tag_350.re;
  assign rcache_line[1][94].status_reg.status = reg2hw.status_350.q;//status_reg_t'(reg2hw.status_350.q);
  assign rcache_line[1][94].status_reg.qe    = reg2hw.status_350.qe;
  assign rcache_line[1][94].status_reg.re    = reg2hw.status_350.re;


  assign rcache_line[1][95].tag_reg.tag      = reg2hw.tag_351.q;
  assign rcache_line[1][95].tag_reg.qe       = reg2hw.tag_351.qe;
  assign rcache_line[1][95].tag_reg.re       = reg2hw.tag_351.re;
  assign rcache_line[1][95].status_reg.status = reg2hw.status_351.q;//status_reg_t'(reg2hw.status_351.q);
  assign rcache_line[1][95].status_reg.qe    = reg2hw.status_351.qe;
  assign rcache_line[1][95].status_reg.re    = reg2hw.status_351.re;


  assign rcache_line[1][96].tag_reg.tag      = reg2hw.tag_352.q;
  assign rcache_line[1][96].tag_reg.qe       = reg2hw.tag_352.qe;
  assign rcache_line[1][96].tag_reg.re       = reg2hw.tag_352.re;
  assign rcache_line[1][96].status_reg.status = reg2hw.status_352.q;//status_reg_t'(reg2hw.status_352.q);
  assign rcache_line[1][96].status_reg.qe    = reg2hw.status_352.qe;
  assign rcache_line[1][96].status_reg.re    = reg2hw.status_352.re;


  assign rcache_line[1][97].tag_reg.tag      = reg2hw.tag_353.q;
  assign rcache_line[1][97].tag_reg.qe       = reg2hw.tag_353.qe;
  assign rcache_line[1][97].tag_reg.re       = reg2hw.tag_353.re;
  assign rcache_line[1][97].status_reg.status = reg2hw.status_353.q;//status_reg_t'(reg2hw.status_353.q);
  assign rcache_line[1][97].status_reg.qe    = reg2hw.status_353.qe;
  assign rcache_line[1][97].status_reg.re    = reg2hw.status_353.re;


  assign rcache_line[1][98].tag_reg.tag      = reg2hw.tag_354.q;
  assign rcache_line[1][98].tag_reg.qe       = reg2hw.tag_354.qe;
  assign rcache_line[1][98].tag_reg.re       = reg2hw.tag_354.re;
  assign rcache_line[1][98].status_reg.status = reg2hw.status_354.q;//status_reg_t'(reg2hw.status_354.q);
  assign rcache_line[1][98].status_reg.qe    = reg2hw.status_354.qe;
  assign rcache_line[1][98].status_reg.re    = reg2hw.status_354.re;


  assign rcache_line[1][99].tag_reg.tag      = reg2hw.tag_355.q;
  assign rcache_line[1][99].tag_reg.qe       = reg2hw.tag_355.qe;
  assign rcache_line[1][99].tag_reg.re       = reg2hw.tag_355.re;
  assign rcache_line[1][99].status_reg.status = reg2hw.status_355.q;//status_reg_t'(reg2hw.status_355.q);
  assign rcache_line[1][99].status_reg.qe    = reg2hw.status_355.qe;
  assign rcache_line[1][99].status_reg.re    = reg2hw.status_355.re;


  assign rcache_line[1][100].tag_reg.tag      = reg2hw.tag_356.q;
  assign rcache_line[1][100].tag_reg.qe       = reg2hw.tag_356.qe;
  assign rcache_line[1][100].tag_reg.re       = reg2hw.tag_356.re;
  assign rcache_line[1][100].status_reg.status = reg2hw.status_356.q;//status_reg_t'(reg2hw.status_356.q);
  assign rcache_line[1][100].status_reg.qe    = reg2hw.status_356.qe;
  assign rcache_line[1][100].status_reg.re    = reg2hw.status_356.re;


  assign rcache_line[1][101].tag_reg.tag      = reg2hw.tag_357.q;
  assign rcache_line[1][101].tag_reg.qe       = reg2hw.tag_357.qe;
  assign rcache_line[1][101].tag_reg.re       = reg2hw.tag_357.re;
  assign rcache_line[1][101].status_reg.status = reg2hw.status_357.q;//status_reg_t'(reg2hw.status_357.q);
  assign rcache_line[1][101].status_reg.qe    = reg2hw.status_357.qe;
  assign rcache_line[1][101].status_reg.re    = reg2hw.status_357.re;


  assign rcache_line[1][102].tag_reg.tag      = reg2hw.tag_358.q;
  assign rcache_line[1][102].tag_reg.qe       = reg2hw.tag_358.qe;
  assign rcache_line[1][102].tag_reg.re       = reg2hw.tag_358.re;
  assign rcache_line[1][102].status_reg.status = reg2hw.status_358.q;//status_reg_t'(reg2hw.status_358.q);
  assign rcache_line[1][102].status_reg.qe    = reg2hw.status_358.qe;
  assign rcache_line[1][102].status_reg.re    = reg2hw.status_358.re;


  assign rcache_line[1][103].tag_reg.tag      = reg2hw.tag_359.q;
  assign rcache_line[1][103].tag_reg.qe       = reg2hw.tag_359.qe;
  assign rcache_line[1][103].tag_reg.re       = reg2hw.tag_359.re;
  assign rcache_line[1][103].status_reg.status = reg2hw.status_359.q;//status_reg_t'(reg2hw.status_359.q);
  assign rcache_line[1][103].status_reg.qe    = reg2hw.status_359.qe;
  assign rcache_line[1][103].status_reg.re    = reg2hw.status_359.re;


  assign rcache_line[1][104].tag_reg.tag      = reg2hw.tag_360.q;
  assign rcache_line[1][104].tag_reg.qe       = reg2hw.tag_360.qe;
  assign rcache_line[1][104].tag_reg.re       = reg2hw.tag_360.re;
  assign rcache_line[1][104].status_reg.status = reg2hw.status_360.q;//status_reg_t'(reg2hw.status_360.q);
  assign rcache_line[1][104].status_reg.qe    = reg2hw.status_360.qe;
  assign rcache_line[1][104].status_reg.re    = reg2hw.status_360.re;


  assign rcache_line[1][105].tag_reg.tag      = reg2hw.tag_361.q;
  assign rcache_line[1][105].tag_reg.qe       = reg2hw.tag_361.qe;
  assign rcache_line[1][105].tag_reg.re       = reg2hw.tag_361.re;
  assign rcache_line[1][105].status_reg.status = reg2hw.status_361.q;//status_reg_t'(reg2hw.status_361.q);
  assign rcache_line[1][105].status_reg.qe    = reg2hw.status_361.qe;
  assign rcache_line[1][105].status_reg.re    = reg2hw.status_361.re;


  assign rcache_line[1][106].tag_reg.tag      = reg2hw.tag_362.q;
  assign rcache_line[1][106].tag_reg.qe       = reg2hw.tag_362.qe;
  assign rcache_line[1][106].tag_reg.re       = reg2hw.tag_362.re;
  assign rcache_line[1][106].status_reg.status = reg2hw.status_362.q;//status_reg_t'(reg2hw.status_362.q);
  assign rcache_line[1][106].status_reg.qe    = reg2hw.status_362.qe;
  assign rcache_line[1][106].status_reg.re    = reg2hw.status_362.re;


  assign rcache_line[1][107].tag_reg.tag      = reg2hw.tag_363.q;
  assign rcache_line[1][107].tag_reg.qe       = reg2hw.tag_363.qe;
  assign rcache_line[1][107].tag_reg.re       = reg2hw.tag_363.re;
  assign rcache_line[1][107].status_reg.status = reg2hw.status_363.q;//status_reg_t'(reg2hw.status_363.q);
  assign rcache_line[1][107].status_reg.qe    = reg2hw.status_363.qe;
  assign rcache_line[1][107].status_reg.re    = reg2hw.status_363.re;


  assign rcache_line[1][108].tag_reg.tag      = reg2hw.tag_364.q;
  assign rcache_line[1][108].tag_reg.qe       = reg2hw.tag_364.qe;
  assign rcache_line[1][108].tag_reg.re       = reg2hw.tag_364.re;
  assign rcache_line[1][108].status_reg.status = reg2hw.status_364.q;//status_reg_t'(reg2hw.status_364.q);
  assign rcache_line[1][108].status_reg.qe    = reg2hw.status_364.qe;
  assign rcache_line[1][108].status_reg.re    = reg2hw.status_364.re;


  assign rcache_line[1][109].tag_reg.tag      = reg2hw.tag_365.q;
  assign rcache_line[1][109].tag_reg.qe       = reg2hw.tag_365.qe;
  assign rcache_line[1][109].tag_reg.re       = reg2hw.tag_365.re;
  assign rcache_line[1][109].status_reg.status = reg2hw.status_365.q;//status_reg_t'(reg2hw.status_365.q);
  assign rcache_line[1][109].status_reg.qe    = reg2hw.status_365.qe;
  assign rcache_line[1][109].status_reg.re    = reg2hw.status_365.re;


  assign rcache_line[1][110].tag_reg.tag      = reg2hw.tag_366.q;
  assign rcache_line[1][110].tag_reg.qe       = reg2hw.tag_366.qe;
  assign rcache_line[1][110].tag_reg.re       = reg2hw.tag_366.re;
  assign rcache_line[1][110].status_reg.status = reg2hw.status_366.q;//status_reg_t'(reg2hw.status_366.q);
  assign rcache_line[1][110].status_reg.qe    = reg2hw.status_366.qe;
  assign rcache_line[1][110].status_reg.re    = reg2hw.status_366.re;


  assign rcache_line[1][111].tag_reg.tag      = reg2hw.tag_367.q;
  assign rcache_line[1][111].tag_reg.qe       = reg2hw.tag_367.qe;
  assign rcache_line[1][111].tag_reg.re       = reg2hw.tag_367.re;
  assign rcache_line[1][111].status_reg.status = reg2hw.status_367.q;//status_reg_t'(reg2hw.status_367.q);
  assign rcache_line[1][111].status_reg.qe    = reg2hw.status_367.qe;
  assign rcache_line[1][111].status_reg.re    = reg2hw.status_367.re;


  assign rcache_line[1][112].tag_reg.tag      = reg2hw.tag_368.q;
  assign rcache_line[1][112].tag_reg.qe       = reg2hw.tag_368.qe;
  assign rcache_line[1][112].tag_reg.re       = reg2hw.tag_368.re;
  assign rcache_line[1][112].status_reg.status = reg2hw.status_368.q;//status_reg_t'(reg2hw.status_368.q);
  assign rcache_line[1][112].status_reg.qe    = reg2hw.status_368.qe;
  assign rcache_line[1][112].status_reg.re    = reg2hw.status_368.re;


  assign rcache_line[1][113].tag_reg.tag      = reg2hw.tag_369.q;
  assign rcache_line[1][113].tag_reg.qe       = reg2hw.tag_369.qe;
  assign rcache_line[1][113].tag_reg.re       = reg2hw.tag_369.re;
  assign rcache_line[1][113].status_reg.status = reg2hw.status_369.q;//status_reg_t'(reg2hw.status_369.q);
  assign rcache_line[1][113].status_reg.qe    = reg2hw.status_369.qe;
  assign rcache_line[1][113].status_reg.re    = reg2hw.status_369.re;


  assign rcache_line[1][114].tag_reg.tag      = reg2hw.tag_370.q;
  assign rcache_line[1][114].tag_reg.qe       = reg2hw.tag_370.qe;
  assign rcache_line[1][114].tag_reg.re       = reg2hw.tag_370.re;
  assign rcache_line[1][114].status_reg.status = reg2hw.status_370.q;//status_reg_t'(reg2hw.status_370.q);
  assign rcache_line[1][114].status_reg.qe    = reg2hw.status_370.qe;
  assign rcache_line[1][114].status_reg.re    = reg2hw.status_370.re;


  assign rcache_line[1][115].tag_reg.tag      = reg2hw.tag_371.q;
  assign rcache_line[1][115].tag_reg.qe       = reg2hw.tag_371.qe;
  assign rcache_line[1][115].tag_reg.re       = reg2hw.tag_371.re;
  assign rcache_line[1][115].status_reg.status = reg2hw.status_371.q;//status_reg_t'(reg2hw.status_371.q);
  assign rcache_line[1][115].status_reg.qe    = reg2hw.status_371.qe;
  assign rcache_line[1][115].status_reg.re    = reg2hw.status_371.re;


  assign rcache_line[1][116].tag_reg.tag      = reg2hw.tag_372.q;
  assign rcache_line[1][116].tag_reg.qe       = reg2hw.tag_372.qe;
  assign rcache_line[1][116].tag_reg.re       = reg2hw.tag_372.re;
  assign rcache_line[1][116].status_reg.status = reg2hw.status_372.q;//status_reg_t'(reg2hw.status_372.q);
  assign rcache_line[1][116].status_reg.qe    = reg2hw.status_372.qe;
  assign rcache_line[1][116].status_reg.re    = reg2hw.status_372.re;


  assign rcache_line[1][117].tag_reg.tag      = reg2hw.tag_373.q;
  assign rcache_line[1][117].tag_reg.qe       = reg2hw.tag_373.qe;
  assign rcache_line[1][117].tag_reg.re       = reg2hw.tag_373.re;
  assign rcache_line[1][117].status_reg.status = reg2hw.status_373.q;//status_reg_t'(reg2hw.status_373.q);
  assign rcache_line[1][117].status_reg.qe    = reg2hw.status_373.qe;
  assign rcache_line[1][117].status_reg.re    = reg2hw.status_373.re;


  assign rcache_line[1][118].tag_reg.tag      = reg2hw.tag_374.q;
  assign rcache_line[1][118].tag_reg.qe       = reg2hw.tag_374.qe;
  assign rcache_line[1][118].tag_reg.re       = reg2hw.tag_374.re;
  assign rcache_line[1][118].status_reg.status = reg2hw.status_374.q;//status_reg_t'(reg2hw.status_374.q);
  assign rcache_line[1][118].status_reg.qe    = reg2hw.status_374.qe;
  assign rcache_line[1][118].status_reg.re    = reg2hw.status_374.re;


  assign rcache_line[1][119].tag_reg.tag      = reg2hw.tag_375.q;
  assign rcache_line[1][119].tag_reg.qe       = reg2hw.tag_375.qe;
  assign rcache_line[1][119].tag_reg.re       = reg2hw.tag_375.re;
  assign rcache_line[1][119].status_reg.status = reg2hw.status_375.q;//status_reg_t'(reg2hw.status_375.q);
  assign rcache_line[1][119].status_reg.qe    = reg2hw.status_375.qe;
  assign rcache_line[1][119].status_reg.re    = reg2hw.status_375.re;


  assign rcache_line[1][120].tag_reg.tag      = reg2hw.tag_376.q;
  assign rcache_line[1][120].tag_reg.qe       = reg2hw.tag_376.qe;
  assign rcache_line[1][120].tag_reg.re       = reg2hw.tag_376.re;
  assign rcache_line[1][120].status_reg.status = reg2hw.status_376.q;//status_reg_t'(reg2hw.status_376.q);
  assign rcache_line[1][120].status_reg.qe    = reg2hw.status_376.qe;
  assign rcache_line[1][120].status_reg.re    = reg2hw.status_376.re;


  assign rcache_line[1][121].tag_reg.tag      = reg2hw.tag_377.q;
  assign rcache_line[1][121].tag_reg.qe       = reg2hw.tag_377.qe;
  assign rcache_line[1][121].tag_reg.re       = reg2hw.tag_377.re;
  assign rcache_line[1][121].status_reg.status = reg2hw.status_377.q;//status_reg_t'(reg2hw.status_377.q);
  assign rcache_line[1][121].status_reg.qe    = reg2hw.status_377.qe;
  assign rcache_line[1][121].status_reg.re    = reg2hw.status_377.re;


  assign rcache_line[1][122].tag_reg.tag      = reg2hw.tag_378.q;
  assign rcache_line[1][122].tag_reg.qe       = reg2hw.tag_378.qe;
  assign rcache_line[1][122].tag_reg.re       = reg2hw.tag_378.re;
  assign rcache_line[1][122].status_reg.status = reg2hw.status_378.q;//status_reg_t'(reg2hw.status_378.q);
  assign rcache_line[1][122].status_reg.qe    = reg2hw.status_378.qe;
  assign rcache_line[1][122].status_reg.re    = reg2hw.status_378.re;


  assign rcache_line[1][123].tag_reg.tag      = reg2hw.tag_379.q;
  assign rcache_line[1][123].tag_reg.qe       = reg2hw.tag_379.qe;
  assign rcache_line[1][123].tag_reg.re       = reg2hw.tag_379.re;
  assign rcache_line[1][123].status_reg.status = reg2hw.status_379.q;//status_reg_t'(reg2hw.status_379.q);
  assign rcache_line[1][123].status_reg.qe    = reg2hw.status_379.qe;
  assign rcache_line[1][123].status_reg.re    = reg2hw.status_379.re;


  assign rcache_line[1][124].tag_reg.tag      = reg2hw.tag_380.q;
  assign rcache_line[1][124].tag_reg.qe       = reg2hw.tag_380.qe;
  assign rcache_line[1][124].tag_reg.re       = reg2hw.tag_380.re;
  assign rcache_line[1][124].status_reg.status = reg2hw.status_380.q;//status_reg_t'(reg2hw.status_380.q);
  assign rcache_line[1][124].status_reg.qe    = reg2hw.status_380.qe;
  assign rcache_line[1][124].status_reg.re    = reg2hw.status_380.re;


  assign rcache_line[1][125].tag_reg.tag      = reg2hw.tag_381.q;
  assign rcache_line[1][125].tag_reg.qe       = reg2hw.tag_381.qe;
  assign rcache_line[1][125].tag_reg.re       = reg2hw.tag_381.re;
  assign rcache_line[1][125].status_reg.status = reg2hw.status_381.q;//status_reg_t'(reg2hw.status_381.q);
  assign rcache_line[1][125].status_reg.qe    = reg2hw.status_381.qe;
  assign rcache_line[1][125].status_reg.re    = reg2hw.status_381.re;


  assign rcache_line[1][126].tag_reg.tag      = reg2hw.tag_382.q;
  assign rcache_line[1][126].tag_reg.qe       = reg2hw.tag_382.qe;
  assign rcache_line[1][126].tag_reg.re       = reg2hw.tag_382.re;
  assign rcache_line[1][126].status_reg.status = reg2hw.status_382.q;//status_reg_t'(reg2hw.status_382.q);
  assign rcache_line[1][126].status_reg.qe    = reg2hw.status_382.qe;
  assign rcache_line[1][126].status_reg.re    = reg2hw.status_382.re;


  assign rcache_line[1][127].tag_reg.tag      = reg2hw.tag_383.q;
  assign rcache_line[1][127].tag_reg.qe       = reg2hw.tag_383.qe;
  assign rcache_line[1][127].tag_reg.re       = reg2hw.tag_383.re;
  assign rcache_line[1][127].status_reg.status = reg2hw.status_383.q;//status_reg_t'(reg2hw.status_383.q);
  assign rcache_line[1][127].status_reg.qe    = reg2hw.status_383.qe;
  assign rcache_line[1][127].status_reg.re    = reg2hw.status_383.re;


  assign rcache_line[1][128].tag_reg.tag      = reg2hw.tag_384.q;
  assign rcache_line[1][128].tag_reg.qe       = reg2hw.tag_384.qe;
  assign rcache_line[1][128].tag_reg.re       = reg2hw.tag_384.re;
  assign rcache_line[1][128].status_reg.status = reg2hw.status_384.q;//status_reg_t'(reg2hw.status_384.q);
  assign rcache_line[1][128].status_reg.qe    = reg2hw.status_384.qe;
  assign rcache_line[1][128].status_reg.re    = reg2hw.status_384.re;


  assign rcache_line[1][129].tag_reg.tag      = reg2hw.tag_385.q;
  assign rcache_line[1][129].tag_reg.qe       = reg2hw.tag_385.qe;
  assign rcache_line[1][129].tag_reg.re       = reg2hw.tag_385.re;
  assign rcache_line[1][129].status_reg.status = reg2hw.status_385.q;//status_reg_t'(reg2hw.status_385.q);
  assign rcache_line[1][129].status_reg.qe    = reg2hw.status_385.qe;
  assign rcache_line[1][129].status_reg.re    = reg2hw.status_385.re;


  assign rcache_line[1][130].tag_reg.tag      = reg2hw.tag_386.q;
  assign rcache_line[1][130].tag_reg.qe       = reg2hw.tag_386.qe;
  assign rcache_line[1][130].tag_reg.re       = reg2hw.tag_386.re;
  assign rcache_line[1][130].status_reg.status = reg2hw.status_386.q;//status_reg_t'(reg2hw.status_386.q);
  assign rcache_line[1][130].status_reg.qe    = reg2hw.status_386.qe;
  assign rcache_line[1][130].status_reg.re    = reg2hw.status_386.re;


  assign rcache_line[1][131].tag_reg.tag      = reg2hw.tag_387.q;
  assign rcache_line[1][131].tag_reg.qe       = reg2hw.tag_387.qe;
  assign rcache_line[1][131].tag_reg.re       = reg2hw.tag_387.re;
  assign rcache_line[1][131].status_reg.status = reg2hw.status_387.q;//status_reg_t'(reg2hw.status_387.q);
  assign rcache_line[1][131].status_reg.qe    = reg2hw.status_387.qe;
  assign rcache_line[1][131].status_reg.re    = reg2hw.status_387.re;


  assign rcache_line[1][132].tag_reg.tag      = reg2hw.tag_388.q;
  assign rcache_line[1][132].tag_reg.qe       = reg2hw.tag_388.qe;
  assign rcache_line[1][132].tag_reg.re       = reg2hw.tag_388.re;
  assign rcache_line[1][132].status_reg.status = reg2hw.status_388.q;//status_reg_t'(reg2hw.status_388.q);
  assign rcache_line[1][132].status_reg.qe    = reg2hw.status_388.qe;
  assign rcache_line[1][132].status_reg.re    = reg2hw.status_388.re;


  assign rcache_line[1][133].tag_reg.tag      = reg2hw.tag_389.q;
  assign rcache_line[1][133].tag_reg.qe       = reg2hw.tag_389.qe;
  assign rcache_line[1][133].tag_reg.re       = reg2hw.tag_389.re;
  assign rcache_line[1][133].status_reg.status = reg2hw.status_389.q;//status_reg_t'(reg2hw.status_389.q);
  assign rcache_line[1][133].status_reg.qe    = reg2hw.status_389.qe;
  assign rcache_line[1][133].status_reg.re    = reg2hw.status_389.re;


  assign rcache_line[1][134].tag_reg.tag      = reg2hw.tag_390.q;
  assign rcache_line[1][134].tag_reg.qe       = reg2hw.tag_390.qe;
  assign rcache_line[1][134].tag_reg.re       = reg2hw.tag_390.re;
  assign rcache_line[1][134].status_reg.status = reg2hw.status_390.q;//status_reg_t'(reg2hw.status_390.q);
  assign rcache_line[1][134].status_reg.qe    = reg2hw.status_390.qe;
  assign rcache_line[1][134].status_reg.re    = reg2hw.status_390.re;


  assign rcache_line[1][135].tag_reg.tag      = reg2hw.tag_391.q;
  assign rcache_line[1][135].tag_reg.qe       = reg2hw.tag_391.qe;
  assign rcache_line[1][135].tag_reg.re       = reg2hw.tag_391.re;
  assign rcache_line[1][135].status_reg.status = reg2hw.status_391.q;//status_reg_t'(reg2hw.status_391.q);
  assign rcache_line[1][135].status_reg.qe    = reg2hw.status_391.qe;
  assign rcache_line[1][135].status_reg.re    = reg2hw.status_391.re;


  assign rcache_line[1][136].tag_reg.tag      = reg2hw.tag_392.q;
  assign rcache_line[1][136].tag_reg.qe       = reg2hw.tag_392.qe;
  assign rcache_line[1][136].tag_reg.re       = reg2hw.tag_392.re;
  assign rcache_line[1][136].status_reg.status = reg2hw.status_392.q;//status_reg_t'(reg2hw.status_392.q);
  assign rcache_line[1][136].status_reg.qe    = reg2hw.status_392.qe;
  assign rcache_line[1][136].status_reg.re    = reg2hw.status_392.re;


  assign rcache_line[1][137].tag_reg.tag      = reg2hw.tag_393.q;
  assign rcache_line[1][137].tag_reg.qe       = reg2hw.tag_393.qe;
  assign rcache_line[1][137].tag_reg.re       = reg2hw.tag_393.re;
  assign rcache_line[1][137].status_reg.status = reg2hw.status_393.q;//status_reg_t'(reg2hw.status_393.q);
  assign rcache_line[1][137].status_reg.qe    = reg2hw.status_393.qe;
  assign rcache_line[1][137].status_reg.re    = reg2hw.status_393.re;


  assign rcache_line[1][138].tag_reg.tag      = reg2hw.tag_394.q;
  assign rcache_line[1][138].tag_reg.qe       = reg2hw.tag_394.qe;
  assign rcache_line[1][138].tag_reg.re       = reg2hw.tag_394.re;
  assign rcache_line[1][138].status_reg.status = reg2hw.status_394.q;//status_reg_t'(reg2hw.status_394.q);
  assign rcache_line[1][138].status_reg.qe    = reg2hw.status_394.qe;
  assign rcache_line[1][138].status_reg.re    = reg2hw.status_394.re;


  assign rcache_line[1][139].tag_reg.tag      = reg2hw.tag_395.q;
  assign rcache_line[1][139].tag_reg.qe       = reg2hw.tag_395.qe;
  assign rcache_line[1][139].tag_reg.re       = reg2hw.tag_395.re;
  assign rcache_line[1][139].status_reg.status = reg2hw.status_395.q;//status_reg_t'(reg2hw.status_395.q);
  assign rcache_line[1][139].status_reg.qe    = reg2hw.status_395.qe;
  assign rcache_line[1][139].status_reg.re    = reg2hw.status_395.re;


  assign rcache_line[1][140].tag_reg.tag      = reg2hw.tag_396.q;
  assign rcache_line[1][140].tag_reg.qe       = reg2hw.tag_396.qe;
  assign rcache_line[1][140].tag_reg.re       = reg2hw.tag_396.re;
  assign rcache_line[1][140].status_reg.status = reg2hw.status_396.q;//status_reg_t'(reg2hw.status_396.q);
  assign rcache_line[1][140].status_reg.qe    = reg2hw.status_396.qe;
  assign rcache_line[1][140].status_reg.re    = reg2hw.status_396.re;


  assign rcache_line[1][141].tag_reg.tag      = reg2hw.tag_397.q;
  assign rcache_line[1][141].tag_reg.qe       = reg2hw.tag_397.qe;
  assign rcache_line[1][141].tag_reg.re       = reg2hw.tag_397.re;
  assign rcache_line[1][141].status_reg.status = reg2hw.status_397.q;//status_reg_t'(reg2hw.status_397.q);
  assign rcache_line[1][141].status_reg.qe    = reg2hw.status_397.qe;
  assign rcache_line[1][141].status_reg.re    = reg2hw.status_397.re;


  assign rcache_line[1][142].tag_reg.tag      = reg2hw.tag_398.q;
  assign rcache_line[1][142].tag_reg.qe       = reg2hw.tag_398.qe;
  assign rcache_line[1][142].tag_reg.re       = reg2hw.tag_398.re;
  assign rcache_line[1][142].status_reg.status = reg2hw.status_398.q;//status_reg_t'(reg2hw.status_398.q);
  assign rcache_line[1][142].status_reg.qe    = reg2hw.status_398.qe;
  assign rcache_line[1][142].status_reg.re    = reg2hw.status_398.re;


  assign rcache_line[1][143].tag_reg.tag      = reg2hw.tag_399.q;
  assign rcache_line[1][143].tag_reg.qe       = reg2hw.tag_399.qe;
  assign rcache_line[1][143].tag_reg.re       = reg2hw.tag_399.re;
  assign rcache_line[1][143].status_reg.status = reg2hw.status_399.q;//status_reg_t'(reg2hw.status_399.q);
  assign rcache_line[1][143].status_reg.qe    = reg2hw.status_399.qe;
  assign rcache_line[1][143].status_reg.re    = reg2hw.status_399.re;


  assign rcache_line[1][144].tag_reg.tag      = reg2hw.tag_400.q;
  assign rcache_line[1][144].tag_reg.qe       = reg2hw.tag_400.qe;
  assign rcache_line[1][144].tag_reg.re       = reg2hw.tag_400.re;
  assign rcache_line[1][144].status_reg.status = reg2hw.status_400.q;//status_reg_t'(reg2hw.status_400.q);
  assign rcache_line[1][144].status_reg.qe    = reg2hw.status_400.qe;
  assign rcache_line[1][144].status_reg.re    = reg2hw.status_400.re;


  assign rcache_line[1][145].tag_reg.tag      = reg2hw.tag_401.q;
  assign rcache_line[1][145].tag_reg.qe       = reg2hw.tag_401.qe;
  assign rcache_line[1][145].tag_reg.re       = reg2hw.tag_401.re;
  assign rcache_line[1][145].status_reg.status = reg2hw.status_401.q;//status_reg_t'(reg2hw.status_401.q);
  assign rcache_line[1][145].status_reg.qe    = reg2hw.status_401.qe;
  assign rcache_line[1][145].status_reg.re    = reg2hw.status_401.re;


  assign rcache_line[1][146].tag_reg.tag      = reg2hw.tag_402.q;
  assign rcache_line[1][146].tag_reg.qe       = reg2hw.tag_402.qe;
  assign rcache_line[1][146].tag_reg.re       = reg2hw.tag_402.re;
  assign rcache_line[1][146].status_reg.status = reg2hw.status_402.q;//status_reg_t'(reg2hw.status_402.q);
  assign rcache_line[1][146].status_reg.qe    = reg2hw.status_402.qe;
  assign rcache_line[1][146].status_reg.re    = reg2hw.status_402.re;


  assign rcache_line[1][147].tag_reg.tag      = reg2hw.tag_403.q;
  assign rcache_line[1][147].tag_reg.qe       = reg2hw.tag_403.qe;
  assign rcache_line[1][147].tag_reg.re       = reg2hw.tag_403.re;
  assign rcache_line[1][147].status_reg.status = reg2hw.status_403.q;//status_reg_t'(reg2hw.status_403.q);
  assign rcache_line[1][147].status_reg.qe    = reg2hw.status_403.qe;
  assign rcache_line[1][147].status_reg.re    = reg2hw.status_403.re;


  assign rcache_line[1][148].tag_reg.tag      = reg2hw.tag_404.q;
  assign rcache_line[1][148].tag_reg.qe       = reg2hw.tag_404.qe;
  assign rcache_line[1][148].tag_reg.re       = reg2hw.tag_404.re;
  assign rcache_line[1][148].status_reg.status = reg2hw.status_404.q;//status_reg_t'(reg2hw.status_404.q);
  assign rcache_line[1][148].status_reg.qe    = reg2hw.status_404.qe;
  assign rcache_line[1][148].status_reg.re    = reg2hw.status_404.re;


  assign rcache_line[1][149].tag_reg.tag      = reg2hw.tag_405.q;
  assign rcache_line[1][149].tag_reg.qe       = reg2hw.tag_405.qe;
  assign rcache_line[1][149].tag_reg.re       = reg2hw.tag_405.re;
  assign rcache_line[1][149].status_reg.status = reg2hw.status_405.q;//status_reg_t'(reg2hw.status_405.q);
  assign rcache_line[1][149].status_reg.qe    = reg2hw.status_405.qe;
  assign rcache_line[1][149].status_reg.re    = reg2hw.status_405.re;


  assign rcache_line[1][150].tag_reg.tag      = reg2hw.tag_406.q;
  assign rcache_line[1][150].tag_reg.qe       = reg2hw.tag_406.qe;
  assign rcache_line[1][150].tag_reg.re       = reg2hw.tag_406.re;
  assign rcache_line[1][150].status_reg.status = reg2hw.status_406.q;//status_reg_t'(reg2hw.status_406.q);
  assign rcache_line[1][150].status_reg.qe    = reg2hw.status_406.qe;
  assign rcache_line[1][150].status_reg.re    = reg2hw.status_406.re;


  assign rcache_line[1][151].tag_reg.tag      = reg2hw.tag_407.q;
  assign rcache_line[1][151].tag_reg.qe       = reg2hw.tag_407.qe;
  assign rcache_line[1][151].tag_reg.re       = reg2hw.tag_407.re;
  assign rcache_line[1][151].status_reg.status = reg2hw.status_407.q;//status_reg_t'(reg2hw.status_407.q);
  assign rcache_line[1][151].status_reg.qe    = reg2hw.status_407.qe;
  assign rcache_line[1][151].status_reg.re    = reg2hw.status_407.re;


  assign rcache_line[1][152].tag_reg.tag      = reg2hw.tag_408.q;
  assign rcache_line[1][152].tag_reg.qe       = reg2hw.tag_408.qe;
  assign rcache_line[1][152].tag_reg.re       = reg2hw.tag_408.re;
  assign rcache_line[1][152].status_reg.status = reg2hw.status_408.q;//status_reg_t'(reg2hw.status_408.q);
  assign rcache_line[1][152].status_reg.qe    = reg2hw.status_408.qe;
  assign rcache_line[1][152].status_reg.re    = reg2hw.status_408.re;


  assign rcache_line[1][153].tag_reg.tag      = reg2hw.tag_409.q;
  assign rcache_line[1][153].tag_reg.qe       = reg2hw.tag_409.qe;
  assign rcache_line[1][153].tag_reg.re       = reg2hw.tag_409.re;
  assign rcache_line[1][153].status_reg.status = reg2hw.status_409.q;//status_reg_t'(reg2hw.status_409.q);
  assign rcache_line[1][153].status_reg.qe    = reg2hw.status_409.qe;
  assign rcache_line[1][153].status_reg.re    = reg2hw.status_409.re;


  assign rcache_line[1][154].tag_reg.tag      = reg2hw.tag_410.q;
  assign rcache_line[1][154].tag_reg.qe       = reg2hw.tag_410.qe;
  assign rcache_line[1][154].tag_reg.re       = reg2hw.tag_410.re;
  assign rcache_line[1][154].status_reg.status = reg2hw.status_410.q;//status_reg_t'(reg2hw.status_410.q);
  assign rcache_line[1][154].status_reg.qe    = reg2hw.status_410.qe;
  assign rcache_line[1][154].status_reg.re    = reg2hw.status_410.re;


  assign rcache_line[1][155].tag_reg.tag      = reg2hw.tag_411.q;
  assign rcache_line[1][155].tag_reg.qe       = reg2hw.tag_411.qe;
  assign rcache_line[1][155].tag_reg.re       = reg2hw.tag_411.re;
  assign rcache_line[1][155].status_reg.status = reg2hw.status_411.q;//status_reg_t'(reg2hw.status_411.q);
  assign rcache_line[1][155].status_reg.qe    = reg2hw.status_411.qe;
  assign rcache_line[1][155].status_reg.re    = reg2hw.status_411.re;


  assign rcache_line[1][156].tag_reg.tag      = reg2hw.tag_412.q;
  assign rcache_line[1][156].tag_reg.qe       = reg2hw.tag_412.qe;
  assign rcache_line[1][156].tag_reg.re       = reg2hw.tag_412.re;
  assign rcache_line[1][156].status_reg.status = reg2hw.status_412.q;//status_reg_t'(reg2hw.status_412.q);
  assign rcache_line[1][156].status_reg.qe    = reg2hw.status_412.qe;
  assign rcache_line[1][156].status_reg.re    = reg2hw.status_412.re;


  assign rcache_line[1][157].tag_reg.tag      = reg2hw.tag_413.q;
  assign rcache_line[1][157].tag_reg.qe       = reg2hw.tag_413.qe;
  assign rcache_line[1][157].tag_reg.re       = reg2hw.tag_413.re;
  assign rcache_line[1][157].status_reg.status = reg2hw.status_413.q;//status_reg_t'(reg2hw.status_413.q);
  assign rcache_line[1][157].status_reg.qe    = reg2hw.status_413.qe;
  assign rcache_line[1][157].status_reg.re    = reg2hw.status_413.re;


  assign rcache_line[1][158].tag_reg.tag      = reg2hw.tag_414.q;
  assign rcache_line[1][158].tag_reg.qe       = reg2hw.tag_414.qe;
  assign rcache_line[1][158].tag_reg.re       = reg2hw.tag_414.re;
  assign rcache_line[1][158].status_reg.status = reg2hw.status_414.q;//status_reg_t'(reg2hw.status_414.q);
  assign rcache_line[1][158].status_reg.qe    = reg2hw.status_414.qe;
  assign rcache_line[1][158].status_reg.re    = reg2hw.status_414.re;


  assign rcache_line[1][159].tag_reg.tag      = reg2hw.tag_415.q;
  assign rcache_line[1][159].tag_reg.qe       = reg2hw.tag_415.qe;
  assign rcache_line[1][159].tag_reg.re       = reg2hw.tag_415.re;
  assign rcache_line[1][159].status_reg.status = reg2hw.status_415.q;//status_reg_t'(reg2hw.status_415.q);
  assign rcache_line[1][159].status_reg.qe    = reg2hw.status_415.qe;
  assign rcache_line[1][159].status_reg.re    = reg2hw.status_415.re;


  assign rcache_line[1][160].tag_reg.tag      = reg2hw.tag_416.q;
  assign rcache_line[1][160].tag_reg.qe       = reg2hw.tag_416.qe;
  assign rcache_line[1][160].tag_reg.re       = reg2hw.tag_416.re;
  assign rcache_line[1][160].status_reg.status = reg2hw.status_416.q;//status_reg_t'(reg2hw.status_416.q);
  assign rcache_line[1][160].status_reg.qe    = reg2hw.status_416.qe;
  assign rcache_line[1][160].status_reg.re    = reg2hw.status_416.re;


  assign rcache_line[1][161].tag_reg.tag      = reg2hw.tag_417.q;
  assign rcache_line[1][161].tag_reg.qe       = reg2hw.tag_417.qe;
  assign rcache_line[1][161].tag_reg.re       = reg2hw.tag_417.re;
  assign rcache_line[1][161].status_reg.status = reg2hw.status_417.q;//status_reg_t'(reg2hw.status_417.q);
  assign rcache_line[1][161].status_reg.qe    = reg2hw.status_417.qe;
  assign rcache_line[1][161].status_reg.re    = reg2hw.status_417.re;


  assign rcache_line[1][162].tag_reg.tag      = reg2hw.tag_418.q;
  assign rcache_line[1][162].tag_reg.qe       = reg2hw.tag_418.qe;
  assign rcache_line[1][162].tag_reg.re       = reg2hw.tag_418.re;
  assign rcache_line[1][162].status_reg.status = reg2hw.status_418.q;//status_reg_t'(reg2hw.status_418.q);
  assign rcache_line[1][162].status_reg.qe    = reg2hw.status_418.qe;
  assign rcache_line[1][162].status_reg.re    = reg2hw.status_418.re;


  assign rcache_line[1][163].tag_reg.tag      = reg2hw.tag_419.q;
  assign rcache_line[1][163].tag_reg.qe       = reg2hw.tag_419.qe;
  assign rcache_line[1][163].tag_reg.re       = reg2hw.tag_419.re;
  assign rcache_line[1][163].status_reg.status = reg2hw.status_419.q;//status_reg_t'(reg2hw.status_419.q);
  assign rcache_line[1][163].status_reg.qe    = reg2hw.status_419.qe;
  assign rcache_line[1][163].status_reg.re    = reg2hw.status_419.re;


  assign rcache_line[1][164].tag_reg.tag      = reg2hw.tag_420.q;
  assign rcache_line[1][164].tag_reg.qe       = reg2hw.tag_420.qe;
  assign rcache_line[1][164].tag_reg.re       = reg2hw.tag_420.re;
  assign rcache_line[1][164].status_reg.status = reg2hw.status_420.q;//status_reg_t'(reg2hw.status_420.q);
  assign rcache_line[1][164].status_reg.qe    = reg2hw.status_420.qe;
  assign rcache_line[1][164].status_reg.re    = reg2hw.status_420.re;


  assign rcache_line[1][165].tag_reg.tag      = reg2hw.tag_421.q;
  assign rcache_line[1][165].tag_reg.qe       = reg2hw.tag_421.qe;
  assign rcache_line[1][165].tag_reg.re       = reg2hw.tag_421.re;
  assign rcache_line[1][165].status_reg.status = reg2hw.status_421.q;//status_reg_t'(reg2hw.status_421.q);
  assign rcache_line[1][165].status_reg.qe    = reg2hw.status_421.qe;
  assign rcache_line[1][165].status_reg.re    = reg2hw.status_421.re;


  assign rcache_line[1][166].tag_reg.tag      = reg2hw.tag_422.q;
  assign rcache_line[1][166].tag_reg.qe       = reg2hw.tag_422.qe;
  assign rcache_line[1][166].tag_reg.re       = reg2hw.tag_422.re;
  assign rcache_line[1][166].status_reg.status = reg2hw.status_422.q;//status_reg_t'(reg2hw.status_422.q);
  assign rcache_line[1][166].status_reg.qe    = reg2hw.status_422.qe;
  assign rcache_line[1][166].status_reg.re    = reg2hw.status_422.re;


  assign rcache_line[1][167].tag_reg.tag      = reg2hw.tag_423.q;
  assign rcache_line[1][167].tag_reg.qe       = reg2hw.tag_423.qe;
  assign rcache_line[1][167].tag_reg.re       = reg2hw.tag_423.re;
  assign rcache_line[1][167].status_reg.status = reg2hw.status_423.q;//status_reg_t'(reg2hw.status_423.q);
  assign rcache_line[1][167].status_reg.qe    = reg2hw.status_423.qe;
  assign rcache_line[1][167].status_reg.re    = reg2hw.status_423.re;


  assign rcache_line[1][168].tag_reg.tag      = reg2hw.tag_424.q;
  assign rcache_line[1][168].tag_reg.qe       = reg2hw.tag_424.qe;
  assign rcache_line[1][168].tag_reg.re       = reg2hw.tag_424.re;
  assign rcache_line[1][168].status_reg.status = reg2hw.status_424.q;//status_reg_t'(reg2hw.status_424.q);
  assign rcache_line[1][168].status_reg.qe    = reg2hw.status_424.qe;
  assign rcache_line[1][168].status_reg.re    = reg2hw.status_424.re;


  assign rcache_line[1][169].tag_reg.tag      = reg2hw.tag_425.q;
  assign rcache_line[1][169].tag_reg.qe       = reg2hw.tag_425.qe;
  assign rcache_line[1][169].tag_reg.re       = reg2hw.tag_425.re;
  assign rcache_line[1][169].status_reg.status = reg2hw.status_425.q;//status_reg_t'(reg2hw.status_425.q);
  assign rcache_line[1][169].status_reg.qe    = reg2hw.status_425.qe;
  assign rcache_line[1][169].status_reg.re    = reg2hw.status_425.re;


  assign rcache_line[1][170].tag_reg.tag      = reg2hw.tag_426.q;
  assign rcache_line[1][170].tag_reg.qe       = reg2hw.tag_426.qe;
  assign rcache_line[1][170].tag_reg.re       = reg2hw.tag_426.re;
  assign rcache_line[1][170].status_reg.status = reg2hw.status_426.q;//status_reg_t'(reg2hw.status_426.q);
  assign rcache_line[1][170].status_reg.qe    = reg2hw.status_426.qe;
  assign rcache_line[1][170].status_reg.re    = reg2hw.status_426.re;


  assign rcache_line[1][171].tag_reg.tag      = reg2hw.tag_427.q;
  assign rcache_line[1][171].tag_reg.qe       = reg2hw.tag_427.qe;
  assign rcache_line[1][171].tag_reg.re       = reg2hw.tag_427.re;
  assign rcache_line[1][171].status_reg.status = reg2hw.status_427.q;//status_reg_t'(reg2hw.status_427.q);
  assign rcache_line[1][171].status_reg.qe    = reg2hw.status_427.qe;
  assign rcache_line[1][171].status_reg.re    = reg2hw.status_427.re;


  assign rcache_line[1][172].tag_reg.tag      = reg2hw.tag_428.q;
  assign rcache_line[1][172].tag_reg.qe       = reg2hw.tag_428.qe;
  assign rcache_line[1][172].tag_reg.re       = reg2hw.tag_428.re;
  assign rcache_line[1][172].status_reg.status = reg2hw.status_428.q;//status_reg_t'(reg2hw.status_428.q);
  assign rcache_line[1][172].status_reg.qe    = reg2hw.status_428.qe;
  assign rcache_line[1][172].status_reg.re    = reg2hw.status_428.re;


  assign rcache_line[1][173].tag_reg.tag      = reg2hw.tag_429.q;
  assign rcache_line[1][173].tag_reg.qe       = reg2hw.tag_429.qe;
  assign rcache_line[1][173].tag_reg.re       = reg2hw.tag_429.re;
  assign rcache_line[1][173].status_reg.status = reg2hw.status_429.q;//status_reg_t'(reg2hw.status_429.q);
  assign rcache_line[1][173].status_reg.qe    = reg2hw.status_429.qe;
  assign rcache_line[1][173].status_reg.re    = reg2hw.status_429.re;


  assign rcache_line[1][174].tag_reg.tag      = reg2hw.tag_430.q;
  assign rcache_line[1][174].tag_reg.qe       = reg2hw.tag_430.qe;
  assign rcache_line[1][174].tag_reg.re       = reg2hw.tag_430.re;
  assign rcache_line[1][174].status_reg.status = reg2hw.status_430.q;//status_reg_t'(reg2hw.status_430.q);
  assign rcache_line[1][174].status_reg.qe    = reg2hw.status_430.qe;
  assign rcache_line[1][174].status_reg.re    = reg2hw.status_430.re;


  assign rcache_line[1][175].tag_reg.tag      = reg2hw.tag_431.q;
  assign rcache_line[1][175].tag_reg.qe       = reg2hw.tag_431.qe;
  assign rcache_line[1][175].tag_reg.re       = reg2hw.tag_431.re;
  assign rcache_line[1][175].status_reg.status = reg2hw.status_431.q;//status_reg_t'(reg2hw.status_431.q);
  assign rcache_line[1][175].status_reg.qe    = reg2hw.status_431.qe;
  assign rcache_line[1][175].status_reg.re    = reg2hw.status_431.re;


  assign rcache_line[1][176].tag_reg.tag      = reg2hw.tag_432.q;
  assign rcache_line[1][176].tag_reg.qe       = reg2hw.tag_432.qe;
  assign rcache_line[1][176].tag_reg.re       = reg2hw.tag_432.re;
  assign rcache_line[1][176].status_reg.status = reg2hw.status_432.q;//status_reg_t'(reg2hw.status_432.q);
  assign rcache_line[1][176].status_reg.qe    = reg2hw.status_432.qe;
  assign rcache_line[1][176].status_reg.re    = reg2hw.status_432.re;


  assign rcache_line[1][177].tag_reg.tag      = reg2hw.tag_433.q;
  assign rcache_line[1][177].tag_reg.qe       = reg2hw.tag_433.qe;
  assign rcache_line[1][177].tag_reg.re       = reg2hw.tag_433.re;
  assign rcache_line[1][177].status_reg.status = reg2hw.status_433.q;//status_reg_t'(reg2hw.status_433.q);
  assign rcache_line[1][177].status_reg.qe    = reg2hw.status_433.qe;
  assign rcache_line[1][177].status_reg.re    = reg2hw.status_433.re;


  assign rcache_line[1][178].tag_reg.tag      = reg2hw.tag_434.q;
  assign rcache_line[1][178].tag_reg.qe       = reg2hw.tag_434.qe;
  assign rcache_line[1][178].tag_reg.re       = reg2hw.tag_434.re;
  assign rcache_line[1][178].status_reg.status = reg2hw.status_434.q;//status_reg_t'(reg2hw.status_434.q);
  assign rcache_line[1][178].status_reg.qe    = reg2hw.status_434.qe;
  assign rcache_line[1][178].status_reg.re    = reg2hw.status_434.re;


  assign rcache_line[1][179].tag_reg.tag      = reg2hw.tag_435.q;
  assign rcache_line[1][179].tag_reg.qe       = reg2hw.tag_435.qe;
  assign rcache_line[1][179].tag_reg.re       = reg2hw.tag_435.re;
  assign rcache_line[1][179].status_reg.status = reg2hw.status_435.q;//status_reg_t'(reg2hw.status_435.q);
  assign rcache_line[1][179].status_reg.qe    = reg2hw.status_435.qe;
  assign rcache_line[1][179].status_reg.re    = reg2hw.status_435.re;


  assign rcache_line[1][180].tag_reg.tag      = reg2hw.tag_436.q;
  assign rcache_line[1][180].tag_reg.qe       = reg2hw.tag_436.qe;
  assign rcache_line[1][180].tag_reg.re       = reg2hw.tag_436.re;
  assign rcache_line[1][180].status_reg.status = reg2hw.status_436.q;//status_reg_t'(reg2hw.status_436.q);
  assign rcache_line[1][180].status_reg.qe    = reg2hw.status_436.qe;
  assign rcache_line[1][180].status_reg.re    = reg2hw.status_436.re;


  assign rcache_line[1][181].tag_reg.tag      = reg2hw.tag_437.q;
  assign rcache_line[1][181].tag_reg.qe       = reg2hw.tag_437.qe;
  assign rcache_line[1][181].tag_reg.re       = reg2hw.tag_437.re;
  assign rcache_line[1][181].status_reg.status = reg2hw.status_437.q;//status_reg_t'(reg2hw.status_437.q);
  assign rcache_line[1][181].status_reg.qe    = reg2hw.status_437.qe;
  assign rcache_line[1][181].status_reg.re    = reg2hw.status_437.re;


  assign rcache_line[1][182].tag_reg.tag      = reg2hw.tag_438.q;
  assign rcache_line[1][182].tag_reg.qe       = reg2hw.tag_438.qe;
  assign rcache_line[1][182].tag_reg.re       = reg2hw.tag_438.re;
  assign rcache_line[1][182].status_reg.status = reg2hw.status_438.q;//status_reg_t'(reg2hw.status_438.q);
  assign rcache_line[1][182].status_reg.qe    = reg2hw.status_438.qe;
  assign rcache_line[1][182].status_reg.re    = reg2hw.status_438.re;


  assign rcache_line[1][183].tag_reg.tag      = reg2hw.tag_439.q;
  assign rcache_line[1][183].tag_reg.qe       = reg2hw.tag_439.qe;
  assign rcache_line[1][183].tag_reg.re       = reg2hw.tag_439.re;
  assign rcache_line[1][183].status_reg.status = reg2hw.status_439.q;//status_reg_t'(reg2hw.status_439.q);
  assign rcache_line[1][183].status_reg.qe    = reg2hw.status_439.qe;
  assign rcache_line[1][183].status_reg.re    = reg2hw.status_439.re;


  assign rcache_line[1][184].tag_reg.tag      = reg2hw.tag_440.q;
  assign rcache_line[1][184].tag_reg.qe       = reg2hw.tag_440.qe;
  assign rcache_line[1][184].tag_reg.re       = reg2hw.tag_440.re;
  assign rcache_line[1][184].status_reg.status = reg2hw.status_440.q;//status_reg_t'(reg2hw.status_440.q);
  assign rcache_line[1][184].status_reg.qe    = reg2hw.status_440.qe;
  assign rcache_line[1][184].status_reg.re    = reg2hw.status_440.re;


  assign rcache_line[1][185].tag_reg.tag      = reg2hw.tag_441.q;
  assign rcache_line[1][185].tag_reg.qe       = reg2hw.tag_441.qe;
  assign rcache_line[1][185].tag_reg.re       = reg2hw.tag_441.re;
  assign rcache_line[1][185].status_reg.status = reg2hw.status_441.q;//status_reg_t'(reg2hw.status_441.q);
  assign rcache_line[1][185].status_reg.qe    = reg2hw.status_441.qe;
  assign rcache_line[1][185].status_reg.re    = reg2hw.status_441.re;


  assign rcache_line[1][186].tag_reg.tag      = reg2hw.tag_442.q;
  assign rcache_line[1][186].tag_reg.qe       = reg2hw.tag_442.qe;
  assign rcache_line[1][186].tag_reg.re       = reg2hw.tag_442.re;
  assign rcache_line[1][186].status_reg.status = reg2hw.status_442.q;//status_reg_t'(reg2hw.status_442.q);
  assign rcache_line[1][186].status_reg.qe    = reg2hw.status_442.qe;
  assign rcache_line[1][186].status_reg.re    = reg2hw.status_442.re;


  assign rcache_line[1][187].tag_reg.tag      = reg2hw.tag_443.q;
  assign rcache_line[1][187].tag_reg.qe       = reg2hw.tag_443.qe;
  assign rcache_line[1][187].tag_reg.re       = reg2hw.tag_443.re;
  assign rcache_line[1][187].status_reg.status = reg2hw.status_443.q;//status_reg_t'(reg2hw.status_443.q);
  assign rcache_line[1][187].status_reg.qe    = reg2hw.status_443.qe;
  assign rcache_line[1][187].status_reg.re    = reg2hw.status_443.re;


  assign rcache_line[1][188].tag_reg.tag      = reg2hw.tag_444.q;
  assign rcache_line[1][188].tag_reg.qe       = reg2hw.tag_444.qe;
  assign rcache_line[1][188].tag_reg.re       = reg2hw.tag_444.re;
  assign rcache_line[1][188].status_reg.status = reg2hw.status_444.q;//status_reg_t'(reg2hw.status_444.q);
  assign rcache_line[1][188].status_reg.qe    = reg2hw.status_444.qe;
  assign rcache_line[1][188].status_reg.re    = reg2hw.status_444.re;


  assign rcache_line[1][189].tag_reg.tag      = reg2hw.tag_445.q;
  assign rcache_line[1][189].tag_reg.qe       = reg2hw.tag_445.qe;
  assign rcache_line[1][189].tag_reg.re       = reg2hw.tag_445.re;
  assign rcache_line[1][189].status_reg.status = reg2hw.status_445.q;//status_reg_t'(reg2hw.status_445.q);
  assign rcache_line[1][189].status_reg.qe    = reg2hw.status_445.qe;
  assign rcache_line[1][189].status_reg.re    = reg2hw.status_445.re;


  assign rcache_line[1][190].tag_reg.tag      = reg2hw.tag_446.q;
  assign rcache_line[1][190].tag_reg.qe       = reg2hw.tag_446.qe;
  assign rcache_line[1][190].tag_reg.re       = reg2hw.tag_446.re;
  assign rcache_line[1][190].status_reg.status = reg2hw.status_446.q;//status_reg_t'(reg2hw.status_446.q);
  assign rcache_line[1][190].status_reg.qe    = reg2hw.status_446.qe;
  assign rcache_line[1][190].status_reg.re    = reg2hw.status_446.re;


  assign rcache_line[1][191].tag_reg.tag      = reg2hw.tag_447.q;
  assign rcache_line[1][191].tag_reg.qe       = reg2hw.tag_447.qe;
  assign rcache_line[1][191].tag_reg.re       = reg2hw.tag_447.re;
  assign rcache_line[1][191].status_reg.status = reg2hw.status_447.q;//status_reg_t'(reg2hw.status_447.q);
  assign rcache_line[1][191].status_reg.qe    = reg2hw.status_447.qe;
  assign rcache_line[1][191].status_reg.re    = reg2hw.status_447.re;


  assign rcache_line[1][192].tag_reg.tag      = reg2hw.tag_448.q;
  assign rcache_line[1][192].tag_reg.qe       = reg2hw.tag_448.qe;
  assign rcache_line[1][192].tag_reg.re       = reg2hw.tag_448.re;
  assign rcache_line[1][192].status_reg.status = reg2hw.status_448.q;//status_reg_t'(reg2hw.status_448.q);
  assign rcache_line[1][192].status_reg.qe    = reg2hw.status_448.qe;
  assign rcache_line[1][192].status_reg.re    = reg2hw.status_448.re;


  assign rcache_line[1][193].tag_reg.tag      = reg2hw.tag_449.q;
  assign rcache_line[1][193].tag_reg.qe       = reg2hw.tag_449.qe;
  assign rcache_line[1][193].tag_reg.re       = reg2hw.tag_449.re;
  assign rcache_line[1][193].status_reg.status = reg2hw.status_449.q;//status_reg_t'(reg2hw.status_449.q);
  assign rcache_line[1][193].status_reg.qe    = reg2hw.status_449.qe;
  assign rcache_line[1][193].status_reg.re    = reg2hw.status_449.re;


  assign rcache_line[1][194].tag_reg.tag      = reg2hw.tag_450.q;
  assign rcache_line[1][194].tag_reg.qe       = reg2hw.tag_450.qe;
  assign rcache_line[1][194].tag_reg.re       = reg2hw.tag_450.re;
  assign rcache_line[1][194].status_reg.status = reg2hw.status_450.q;//status_reg_t'(reg2hw.status_450.q);
  assign rcache_line[1][194].status_reg.qe    = reg2hw.status_450.qe;
  assign rcache_line[1][194].status_reg.re    = reg2hw.status_450.re;


  assign rcache_line[1][195].tag_reg.tag      = reg2hw.tag_451.q;
  assign rcache_line[1][195].tag_reg.qe       = reg2hw.tag_451.qe;
  assign rcache_line[1][195].tag_reg.re       = reg2hw.tag_451.re;
  assign rcache_line[1][195].status_reg.status = reg2hw.status_451.q;//status_reg_t'(reg2hw.status_451.q);
  assign rcache_line[1][195].status_reg.qe    = reg2hw.status_451.qe;
  assign rcache_line[1][195].status_reg.re    = reg2hw.status_451.re;


  assign rcache_line[1][196].tag_reg.tag      = reg2hw.tag_452.q;
  assign rcache_line[1][196].tag_reg.qe       = reg2hw.tag_452.qe;
  assign rcache_line[1][196].tag_reg.re       = reg2hw.tag_452.re;
  assign rcache_line[1][196].status_reg.status = reg2hw.status_452.q;//status_reg_t'(reg2hw.status_452.q);
  assign rcache_line[1][196].status_reg.qe    = reg2hw.status_452.qe;
  assign rcache_line[1][196].status_reg.re    = reg2hw.status_452.re;


  assign rcache_line[1][197].tag_reg.tag      = reg2hw.tag_453.q;
  assign rcache_line[1][197].tag_reg.qe       = reg2hw.tag_453.qe;
  assign rcache_line[1][197].tag_reg.re       = reg2hw.tag_453.re;
  assign rcache_line[1][197].status_reg.status = reg2hw.status_453.q;//status_reg_t'(reg2hw.status_453.q);
  assign rcache_line[1][197].status_reg.qe    = reg2hw.status_453.qe;
  assign rcache_line[1][197].status_reg.re    = reg2hw.status_453.re;


  assign rcache_line[1][198].tag_reg.tag      = reg2hw.tag_454.q;
  assign rcache_line[1][198].tag_reg.qe       = reg2hw.tag_454.qe;
  assign rcache_line[1][198].tag_reg.re       = reg2hw.tag_454.re;
  assign rcache_line[1][198].status_reg.status = reg2hw.status_454.q;//status_reg_t'(reg2hw.status_454.q);
  assign rcache_line[1][198].status_reg.qe    = reg2hw.status_454.qe;
  assign rcache_line[1][198].status_reg.re    = reg2hw.status_454.re;


  assign rcache_line[1][199].tag_reg.tag      = reg2hw.tag_455.q;
  assign rcache_line[1][199].tag_reg.qe       = reg2hw.tag_455.qe;
  assign rcache_line[1][199].tag_reg.re       = reg2hw.tag_455.re;
  assign rcache_line[1][199].status_reg.status = reg2hw.status_455.q;//status_reg_t'(reg2hw.status_455.q);
  assign rcache_line[1][199].status_reg.qe    = reg2hw.status_455.qe;
  assign rcache_line[1][199].status_reg.re    = reg2hw.status_455.re;


  assign rcache_line[1][200].tag_reg.tag      = reg2hw.tag_456.q;
  assign rcache_line[1][200].tag_reg.qe       = reg2hw.tag_456.qe;
  assign rcache_line[1][200].tag_reg.re       = reg2hw.tag_456.re;
  assign rcache_line[1][200].status_reg.status = reg2hw.status_456.q;//status_reg_t'(reg2hw.status_456.q);
  assign rcache_line[1][200].status_reg.qe    = reg2hw.status_456.qe;
  assign rcache_line[1][200].status_reg.re    = reg2hw.status_456.re;


  assign rcache_line[1][201].tag_reg.tag      = reg2hw.tag_457.q;
  assign rcache_line[1][201].tag_reg.qe       = reg2hw.tag_457.qe;
  assign rcache_line[1][201].tag_reg.re       = reg2hw.tag_457.re;
  assign rcache_line[1][201].status_reg.status = reg2hw.status_457.q;//status_reg_t'(reg2hw.status_457.q);
  assign rcache_line[1][201].status_reg.qe    = reg2hw.status_457.qe;
  assign rcache_line[1][201].status_reg.re    = reg2hw.status_457.re;


  assign rcache_line[1][202].tag_reg.tag      = reg2hw.tag_458.q;
  assign rcache_line[1][202].tag_reg.qe       = reg2hw.tag_458.qe;
  assign rcache_line[1][202].tag_reg.re       = reg2hw.tag_458.re;
  assign rcache_line[1][202].status_reg.status = reg2hw.status_458.q;//status_reg_t'(reg2hw.status_458.q);
  assign rcache_line[1][202].status_reg.qe    = reg2hw.status_458.qe;
  assign rcache_line[1][202].status_reg.re    = reg2hw.status_458.re;


  assign rcache_line[1][203].tag_reg.tag      = reg2hw.tag_459.q;
  assign rcache_line[1][203].tag_reg.qe       = reg2hw.tag_459.qe;
  assign rcache_line[1][203].tag_reg.re       = reg2hw.tag_459.re;
  assign rcache_line[1][203].status_reg.status = reg2hw.status_459.q;//status_reg_t'(reg2hw.status_459.q);
  assign rcache_line[1][203].status_reg.qe    = reg2hw.status_459.qe;
  assign rcache_line[1][203].status_reg.re    = reg2hw.status_459.re;


  assign rcache_line[1][204].tag_reg.tag      = reg2hw.tag_460.q;
  assign rcache_line[1][204].tag_reg.qe       = reg2hw.tag_460.qe;
  assign rcache_line[1][204].tag_reg.re       = reg2hw.tag_460.re;
  assign rcache_line[1][204].status_reg.status = reg2hw.status_460.q;//status_reg_t'(reg2hw.status_460.q);
  assign rcache_line[1][204].status_reg.qe    = reg2hw.status_460.qe;
  assign rcache_line[1][204].status_reg.re    = reg2hw.status_460.re;


  assign rcache_line[1][205].tag_reg.tag      = reg2hw.tag_461.q;
  assign rcache_line[1][205].tag_reg.qe       = reg2hw.tag_461.qe;
  assign rcache_line[1][205].tag_reg.re       = reg2hw.tag_461.re;
  assign rcache_line[1][205].status_reg.status = reg2hw.status_461.q;//status_reg_t'(reg2hw.status_461.q);
  assign rcache_line[1][205].status_reg.qe    = reg2hw.status_461.qe;
  assign rcache_line[1][205].status_reg.re    = reg2hw.status_461.re;


  assign rcache_line[1][206].tag_reg.tag      = reg2hw.tag_462.q;
  assign rcache_line[1][206].tag_reg.qe       = reg2hw.tag_462.qe;
  assign rcache_line[1][206].tag_reg.re       = reg2hw.tag_462.re;
  assign rcache_line[1][206].status_reg.status = reg2hw.status_462.q;//status_reg_t'(reg2hw.status_462.q);
  assign rcache_line[1][206].status_reg.qe    = reg2hw.status_462.qe;
  assign rcache_line[1][206].status_reg.re    = reg2hw.status_462.re;


  assign rcache_line[1][207].tag_reg.tag      = reg2hw.tag_463.q;
  assign rcache_line[1][207].tag_reg.qe       = reg2hw.tag_463.qe;
  assign rcache_line[1][207].tag_reg.re       = reg2hw.tag_463.re;
  assign rcache_line[1][207].status_reg.status = reg2hw.status_463.q;//status_reg_t'(reg2hw.status_463.q);
  assign rcache_line[1][207].status_reg.qe    = reg2hw.status_463.qe;
  assign rcache_line[1][207].status_reg.re    = reg2hw.status_463.re;


  assign rcache_line[1][208].tag_reg.tag      = reg2hw.tag_464.q;
  assign rcache_line[1][208].tag_reg.qe       = reg2hw.tag_464.qe;
  assign rcache_line[1][208].tag_reg.re       = reg2hw.tag_464.re;
  assign rcache_line[1][208].status_reg.status = reg2hw.status_464.q;//status_reg_t'(reg2hw.status_464.q);
  assign rcache_line[1][208].status_reg.qe    = reg2hw.status_464.qe;
  assign rcache_line[1][208].status_reg.re    = reg2hw.status_464.re;


  assign rcache_line[1][209].tag_reg.tag      = reg2hw.tag_465.q;
  assign rcache_line[1][209].tag_reg.qe       = reg2hw.tag_465.qe;
  assign rcache_line[1][209].tag_reg.re       = reg2hw.tag_465.re;
  assign rcache_line[1][209].status_reg.status = reg2hw.status_465.q;//status_reg_t'(reg2hw.status_465.q);
  assign rcache_line[1][209].status_reg.qe    = reg2hw.status_465.qe;
  assign rcache_line[1][209].status_reg.re    = reg2hw.status_465.re;


  assign rcache_line[1][210].tag_reg.tag      = reg2hw.tag_466.q;
  assign rcache_line[1][210].tag_reg.qe       = reg2hw.tag_466.qe;
  assign rcache_line[1][210].tag_reg.re       = reg2hw.tag_466.re;
  assign rcache_line[1][210].status_reg.status = reg2hw.status_466.q;//status_reg_t'(reg2hw.status_466.q);
  assign rcache_line[1][210].status_reg.qe    = reg2hw.status_466.qe;
  assign rcache_line[1][210].status_reg.re    = reg2hw.status_466.re;


  assign rcache_line[1][211].tag_reg.tag      = reg2hw.tag_467.q;
  assign rcache_line[1][211].tag_reg.qe       = reg2hw.tag_467.qe;
  assign rcache_line[1][211].tag_reg.re       = reg2hw.tag_467.re;
  assign rcache_line[1][211].status_reg.status = reg2hw.status_467.q;//status_reg_t'(reg2hw.status_467.q);
  assign rcache_line[1][211].status_reg.qe    = reg2hw.status_467.qe;
  assign rcache_line[1][211].status_reg.re    = reg2hw.status_467.re;


  assign rcache_line[1][212].tag_reg.tag      = reg2hw.tag_468.q;
  assign rcache_line[1][212].tag_reg.qe       = reg2hw.tag_468.qe;
  assign rcache_line[1][212].tag_reg.re       = reg2hw.tag_468.re;
  assign rcache_line[1][212].status_reg.status = reg2hw.status_468.q;//status_reg_t'(reg2hw.status_468.q);
  assign rcache_line[1][212].status_reg.qe    = reg2hw.status_468.qe;
  assign rcache_line[1][212].status_reg.re    = reg2hw.status_468.re;


  assign rcache_line[1][213].tag_reg.tag      = reg2hw.tag_469.q;
  assign rcache_line[1][213].tag_reg.qe       = reg2hw.tag_469.qe;
  assign rcache_line[1][213].tag_reg.re       = reg2hw.tag_469.re;
  assign rcache_line[1][213].status_reg.status = reg2hw.status_469.q;//status_reg_t'(reg2hw.status_469.q);
  assign rcache_line[1][213].status_reg.qe    = reg2hw.status_469.qe;
  assign rcache_line[1][213].status_reg.re    = reg2hw.status_469.re;


  assign rcache_line[1][214].tag_reg.tag      = reg2hw.tag_470.q;
  assign rcache_line[1][214].tag_reg.qe       = reg2hw.tag_470.qe;
  assign rcache_line[1][214].tag_reg.re       = reg2hw.tag_470.re;
  assign rcache_line[1][214].status_reg.status = reg2hw.status_470.q;//status_reg_t'(reg2hw.status_470.q);
  assign rcache_line[1][214].status_reg.qe    = reg2hw.status_470.qe;
  assign rcache_line[1][214].status_reg.re    = reg2hw.status_470.re;


  assign rcache_line[1][215].tag_reg.tag      = reg2hw.tag_471.q;
  assign rcache_line[1][215].tag_reg.qe       = reg2hw.tag_471.qe;
  assign rcache_line[1][215].tag_reg.re       = reg2hw.tag_471.re;
  assign rcache_line[1][215].status_reg.status = reg2hw.status_471.q;//status_reg_t'(reg2hw.status_471.q);
  assign rcache_line[1][215].status_reg.qe    = reg2hw.status_471.qe;
  assign rcache_line[1][215].status_reg.re    = reg2hw.status_471.re;


  assign rcache_line[1][216].tag_reg.tag      = reg2hw.tag_472.q;
  assign rcache_line[1][216].tag_reg.qe       = reg2hw.tag_472.qe;
  assign rcache_line[1][216].tag_reg.re       = reg2hw.tag_472.re;
  assign rcache_line[1][216].status_reg.status = reg2hw.status_472.q;//status_reg_t'(reg2hw.status_472.q);
  assign rcache_line[1][216].status_reg.qe    = reg2hw.status_472.qe;
  assign rcache_line[1][216].status_reg.re    = reg2hw.status_472.re;


  assign rcache_line[1][217].tag_reg.tag      = reg2hw.tag_473.q;
  assign rcache_line[1][217].tag_reg.qe       = reg2hw.tag_473.qe;
  assign rcache_line[1][217].tag_reg.re       = reg2hw.tag_473.re;
  assign rcache_line[1][217].status_reg.status = reg2hw.status_473.q;//status_reg_t'(reg2hw.status_473.q);
  assign rcache_line[1][217].status_reg.qe    = reg2hw.status_473.qe;
  assign rcache_line[1][217].status_reg.re    = reg2hw.status_473.re;


  assign rcache_line[1][218].tag_reg.tag      = reg2hw.tag_474.q;
  assign rcache_line[1][218].tag_reg.qe       = reg2hw.tag_474.qe;
  assign rcache_line[1][218].tag_reg.re       = reg2hw.tag_474.re;
  assign rcache_line[1][218].status_reg.status = reg2hw.status_474.q;//status_reg_t'(reg2hw.status_474.q);
  assign rcache_line[1][218].status_reg.qe    = reg2hw.status_474.qe;
  assign rcache_line[1][218].status_reg.re    = reg2hw.status_474.re;


  assign rcache_line[1][219].tag_reg.tag      = reg2hw.tag_475.q;
  assign rcache_line[1][219].tag_reg.qe       = reg2hw.tag_475.qe;
  assign rcache_line[1][219].tag_reg.re       = reg2hw.tag_475.re;
  assign rcache_line[1][219].status_reg.status = reg2hw.status_475.q;//status_reg_t'(reg2hw.status_475.q);
  assign rcache_line[1][219].status_reg.qe    = reg2hw.status_475.qe;
  assign rcache_line[1][219].status_reg.re    = reg2hw.status_475.re;


  assign rcache_line[1][220].tag_reg.tag      = reg2hw.tag_476.q;
  assign rcache_line[1][220].tag_reg.qe       = reg2hw.tag_476.qe;
  assign rcache_line[1][220].tag_reg.re       = reg2hw.tag_476.re;
  assign rcache_line[1][220].status_reg.status = reg2hw.status_476.q;//status_reg_t'(reg2hw.status_476.q);
  assign rcache_line[1][220].status_reg.qe    = reg2hw.status_476.qe;
  assign rcache_line[1][220].status_reg.re    = reg2hw.status_476.re;


  assign rcache_line[1][221].tag_reg.tag      = reg2hw.tag_477.q;
  assign rcache_line[1][221].tag_reg.qe       = reg2hw.tag_477.qe;
  assign rcache_line[1][221].tag_reg.re       = reg2hw.tag_477.re;
  assign rcache_line[1][221].status_reg.status = reg2hw.status_477.q;//status_reg_t'(reg2hw.status_477.q);
  assign rcache_line[1][221].status_reg.qe    = reg2hw.status_477.qe;
  assign rcache_line[1][221].status_reg.re    = reg2hw.status_477.re;


  assign rcache_line[1][222].tag_reg.tag      = reg2hw.tag_478.q;
  assign rcache_line[1][222].tag_reg.qe       = reg2hw.tag_478.qe;
  assign rcache_line[1][222].tag_reg.re       = reg2hw.tag_478.re;
  assign rcache_line[1][222].status_reg.status = reg2hw.status_478.q;//status_reg_t'(reg2hw.status_478.q);
  assign rcache_line[1][222].status_reg.qe    = reg2hw.status_478.qe;
  assign rcache_line[1][222].status_reg.re    = reg2hw.status_478.re;


  assign rcache_line[1][223].tag_reg.tag      = reg2hw.tag_479.q;
  assign rcache_line[1][223].tag_reg.qe       = reg2hw.tag_479.qe;
  assign rcache_line[1][223].tag_reg.re       = reg2hw.tag_479.re;
  assign rcache_line[1][223].status_reg.status = reg2hw.status_479.q;//status_reg_t'(reg2hw.status_479.q);
  assign rcache_line[1][223].status_reg.qe    = reg2hw.status_479.qe;
  assign rcache_line[1][223].status_reg.re    = reg2hw.status_479.re;


  assign rcache_line[1][224].tag_reg.tag      = reg2hw.tag_480.q;
  assign rcache_line[1][224].tag_reg.qe       = reg2hw.tag_480.qe;
  assign rcache_line[1][224].tag_reg.re       = reg2hw.tag_480.re;
  assign rcache_line[1][224].status_reg.status = reg2hw.status_480.q;//status_reg_t'(reg2hw.status_480.q);
  assign rcache_line[1][224].status_reg.qe    = reg2hw.status_480.qe;
  assign rcache_line[1][224].status_reg.re    = reg2hw.status_480.re;


  assign rcache_line[1][225].tag_reg.tag      = reg2hw.tag_481.q;
  assign rcache_line[1][225].tag_reg.qe       = reg2hw.tag_481.qe;
  assign rcache_line[1][225].tag_reg.re       = reg2hw.tag_481.re;
  assign rcache_line[1][225].status_reg.status = reg2hw.status_481.q;//status_reg_t'(reg2hw.status_481.q);
  assign rcache_line[1][225].status_reg.qe    = reg2hw.status_481.qe;
  assign rcache_line[1][225].status_reg.re    = reg2hw.status_481.re;


  assign rcache_line[1][226].tag_reg.tag      = reg2hw.tag_482.q;
  assign rcache_line[1][226].tag_reg.qe       = reg2hw.tag_482.qe;
  assign rcache_line[1][226].tag_reg.re       = reg2hw.tag_482.re;
  assign rcache_line[1][226].status_reg.status = reg2hw.status_482.q;//status_reg_t'(reg2hw.status_482.q);
  assign rcache_line[1][226].status_reg.qe    = reg2hw.status_482.qe;
  assign rcache_line[1][226].status_reg.re    = reg2hw.status_482.re;


  assign rcache_line[1][227].tag_reg.tag      = reg2hw.tag_483.q;
  assign rcache_line[1][227].tag_reg.qe       = reg2hw.tag_483.qe;
  assign rcache_line[1][227].tag_reg.re       = reg2hw.tag_483.re;
  assign rcache_line[1][227].status_reg.status = reg2hw.status_483.q;//status_reg_t'(reg2hw.status_483.q);
  assign rcache_line[1][227].status_reg.qe    = reg2hw.status_483.qe;
  assign rcache_line[1][227].status_reg.re    = reg2hw.status_483.re;


  assign rcache_line[1][228].tag_reg.tag      = reg2hw.tag_484.q;
  assign rcache_line[1][228].tag_reg.qe       = reg2hw.tag_484.qe;
  assign rcache_line[1][228].tag_reg.re       = reg2hw.tag_484.re;
  assign rcache_line[1][228].status_reg.status = reg2hw.status_484.q;//status_reg_t'(reg2hw.status_484.q);
  assign rcache_line[1][228].status_reg.qe    = reg2hw.status_484.qe;
  assign rcache_line[1][228].status_reg.re    = reg2hw.status_484.re;


  assign rcache_line[1][229].tag_reg.tag      = reg2hw.tag_485.q;
  assign rcache_line[1][229].tag_reg.qe       = reg2hw.tag_485.qe;
  assign rcache_line[1][229].tag_reg.re       = reg2hw.tag_485.re;
  assign rcache_line[1][229].status_reg.status = reg2hw.status_485.q;//status_reg_t'(reg2hw.status_485.q);
  assign rcache_line[1][229].status_reg.qe    = reg2hw.status_485.qe;
  assign rcache_line[1][229].status_reg.re    = reg2hw.status_485.re;


  assign rcache_line[1][230].tag_reg.tag      = reg2hw.tag_486.q;
  assign rcache_line[1][230].tag_reg.qe       = reg2hw.tag_486.qe;
  assign rcache_line[1][230].tag_reg.re       = reg2hw.tag_486.re;
  assign rcache_line[1][230].status_reg.status = reg2hw.status_486.q;//status_reg_t'(reg2hw.status_486.q);
  assign rcache_line[1][230].status_reg.qe    = reg2hw.status_486.qe;
  assign rcache_line[1][230].status_reg.re    = reg2hw.status_486.re;


  assign rcache_line[1][231].tag_reg.tag      = reg2hw.tag_487.q;
  assign rcache_line[1][231].tag_reg.qe       = reg2hw.tag_487.qe;
  assign rcache_line[1][231].tag_reg.re       = reg2hw.tag_487.re;
  assign rcache_line[1][231].status_reg.status = reg2hw.status_487.q;//status_reg_t'(reg2hw.status_487.q);
  assign rcache_line[1][231].status_reg.qe    = reg2hw.status_487.qe;
  assign rcache_line[1][231].status_reg.re    = reg2hw.status_487.re;


  assign rcache_line[1][232].tag_reg.tag      = reg2hw.tag_488.q;
  assign rcache_line[1][232].tag_reg.qe       = reg2hw.tag_488.qe;
  assign rcache_line[1][232].tag_reg.re       = reg2hw.tag_488.re;
  assign rcache_line[1][232].status_reg.status = reg2hw.status_488.q;//status_reg_t'(reg2hw.status_488.q);
  assign rcache_line[1][232].status_reg.qe    = reg2hw.status_488.qe;
  assign rcache_line[1][232].status_reg.re    = reg2hw.status_488.re;


  assign rcache_line[1][233].tag_reg.tag      = reg2hw.tag_489.q;
  assign rcache_line[1][233].tag_reg.qe       = reg2hw.tag_489.qe;
  assign rcache_line[1][233].tag_reg.re       = reg2hw.tag_489.re;
  assign rcache_line[1][233].status_reg.status = reg2hw.status_489.q;//status_reg_t'(reg2hw.status_489.q);
  assign rcache_line[1][233].status_reg.qe    = reg2hw.status_489.qe;
  assign rcache_line[1][233].status_reg.re    = reg2hw.status_489.re;


  assign rcache_line[1][234].tag_reg.tag      = reg2hw.tag_490.q;
  assign rcache_line[1][234].tag_reg.qe       = reg2hw.tag_490.qe;
  assign rcache_line[1][234].tag_reg.re       = reg2hw.tag_490.re;
  assign rcache_line[1][234].status_reg.status = reg2hw.status_490.q;//status_reg_t'(reg2hw.status_490.q);
  assign rcache_line[1][234].status_reg.qe    = reg2hw.status_490.qe;
  assign rcache_line[1][234].status_reg.re    = reg2hw.status_490.re;


  assign rcache_line[1][235].tag_reg.tag      = reg2hw.tag_491.q;
  assign rcache_line[1][235].tag_reg.qe       = reg2hw.tag_491.qe;
  assign rcache_line[1][235].tag_reg.re       = reg2hw.tag_491.re;
  assign rcache_line[1][235].status_reg.status = reg2hw.status_491.q;//status_reg_t'(reg2hw.status_491.q);
  assign rcache_line[1][235].status_reg.qe    = reg2hw.status_491.qe;
  assign rcache_line[1][235].status_reg.re    = reg2hw.status_491.re;


  assign rcache_line[1][236].tag_reg.tag      = reg2hw.tag_492.q;
  assign rcache_line[1][236].tag_reg.qe       = reg2hw.tag_492.qe;
  assign rcache_line[1][236].tag_reg.re       = reg2hw.tag_492.re;
  assign rcache_line[1][236].status_reg.status = reg2hw.status_492.q;//status_reg_t'(reg2hw.status_492.q);
  assign rcache_line[1][236].status_reg.qe    = reg2hw.status_492.qe;
  assign rcache_line[1][236].status_reg.re    = reg2hw.status_492.re;


  assign rcache_line[1][237].tag_reg.tag      = reg2hw.tag_493.q;
  assign rcache_line[1][237].tag_reg.qe       = reg2hw.tag_493.qe;
  assign rcache_line[1][237].tag_reg.re       = reg2hw.tag_493.re;
  assign rcache_line[1][237].status_reg.status = reg2hw.status_493.q;//status_reg_t'(reg2hw.status_493.q);
  assign rcache_line[1][237].status_reg.qe    = reg2hw.status_493.qe;
  assign rcache_line[1][237].status_reg.re    = reg2hw.status_493.re;


  assign rcache_line[1][238].tag_reg.tag      = reg2hw.tag_494.q;
  assign rcache_line[1][238].tag_reg.qe       = reg2hw.tag_494.qe;
  assign rcache_line[1][238].tag_reg.re       = reg2hw.tag_494.re;
  assign rcache_line[1][238].status_reg.status = reg2hw.status_494.q;//status_reg_t'(reg2hw.status_494.q);
  assign rcache_line[1][238].status_reg.qe    = reg2hw.status_494.qe;
  assign rcache_line[1][238].status_reg.re    = reg2hw.status_494.re;


  assign rcache_line[1][239].tag_reg.tag      = reg2hw.tag_495.q;
  assign rcache_line[1][239].tag_reg.qe       = reg2hw.tag_495.qe;
  assign rcache_line[1][239].tag_reg.re       = reg2hw.tag_495.re;
  assign rcache_line[1][239].status_reg.status = reg2hw.status_495.q;//status_reg_t'(reg2hw.status_495.q);
  assign rcache_line[1][239].status_reg.qe    = reg2hw.status_495.qe;
  assign rcache_line[1][239].status_reg.re    = reg2hw.status_495.re;


  assign rcache_line[1][240].tag_reg.tag      = reg2hw.tag_496.q;
  assign rcache_line[1][240].tag_reg.qe       = reg2hw.tag_496.qe;
  assign rcache_line[1][240].tag_reg.re       = reg2hw.tag_496.re;
  assign rcache_line[1][240].status_reg.status = reg2hw.status_496.q;//status_reg_t'(reg2hw.status_496.q);
  assign rcache_line[1][240].status_reg.qe    = reg2hw.status_496.qe;
  assign rcache_line[1][240].status_reg.re    = reg2hw.status_496.re;


  assign rcache_line[1][241].tag_reg.tag      = reg2hw.tag_497.q;
  assign rcache_line[1][241].tag_reg.qe       = reg2hw.tag_497.qe;
  assign rcache_line[1][241].tag_reg.re       = reg2hw.tag_497.re;
  assign rcache_line[1][241].status_reg.status = reg2hw.status_497.q;//status_reg_t'(reg2hw.status_497.q);
  assign rcache_line[1][241].status_reg.qe    = reg2hw.status_497.qe;
  assign rcache_line[1][241].status_reg.re    = reg2hw.status_497.re;


  assign rcache_line[1][242].tag_reg.tag      = reg2hw.tag_498.q;
  assign rcache_line[1][242].tag_reg.qe       = reg2hw.tag_498.qe;
  assign rcache_line[1][242].tag_reg.re       = reg2hw.tag_498.re;
  assign rcache_line[1][242].status_reg.status = reg2hw.status_498.q;//status_reg_t'(reg2hw.status_498.q);
  assign rcache_line[1][242].status_reg.qe    = reg2hw.status_498.qe;
  assign rcache_line[1][242].status_reg.re    = reg2hw.status_498.re;


  assign rcache_line[1][243].tag_reg.tag      = reg2hw.tag_499.q;
  assign rcache_line[1][243].tag_reg.qe       = reg2hw.tag_499.qe;
  assign rcache_line[1][243].tag_reg.re       = reg2hw.tag_499.re;
  assign rcache_line[1][243].status_reg.status = reg2hw.status_499.q;//status_reg_t'(reg2hw.status_499.q);
  assign rcache_line[1][243].status_reg.qe    = reg2hw.status_499.qe;
  assign rcache_line[1][243].status_reg.re    = reg2hw.status_499.re;


  assign rcache_line[1][244].tag_reg.tag      = reg2hw.tag_500.q;
  assign rcache_line[1][244].tag_reg.qe       = reg2hw.tag_500.qe;
  assign rcache_line[1][244].tag_reg.re       = reg2hw.tag_500.re;
  assign rcache_line[1][244].status_reg.status = reg2hw.status_500.q;//status_reg_t'(reg2hw.status_500.q);
  assign rcache_line[1][244].status_reg.qe    = reg2hw.status_500.qe;
  assign rcache_line[1][244].status_reg.re    = reg2hw.status_500.re;


  assign rcache_line[1][245].tag_reg.tag      = reg2hw.tag_501.q;
  assign rcache_line[1][245].tag_reg.qe       = reg2hw.tag_501.qe;
  assign rcache_line[1][245].tag_reg.re       = reg2hw.tag_501.re;
  assign rcache_line[1][245].status_reg.status = reg2hw.status_501.q;//status_reg_t'(reg2hw.status_501.q);
  assign rcache_line[1][245].status_reg.qe    = reg2hw.status_501.qe;
  assign rcache_line[1][245].status_reg.re    = reg2hw.status_501.re;


  assign rcache_line[1][246].tag_reg.tag      = reg2hw.tag_502.q;
  assign rcache_line[1][246].tag_reg.qe       = reg2hw.tag_502.qe;
  assign rcache_line[1][246].tag_reg.re       = reg2hw.tag_502.re;
  assign rcache_line[1][246].status_reg.status = reg2hw.status_502.q;//status_reg_t'(reg2hw.status_502.q);
  assign rcache_line[1][246].status_reg.qe    = reg2hw.status_502.qe;
  assign rcache_line[1][246].status_reg.re    = reg2hw.status_502.re;


  assign rcache_line[1][247].tag_reg.tag      = reg2hw.tag_503.q;
  assign rcache_line[1][247].tag_reg.qe       = reg2hw.tag_503.qe;
  assign rcache_line[1][247].tag_reg.re       = reg2hw.tag_503.re;
  assign rcache_line[1][247].status_reg.status = reg2hw.status_503.q;//status_reg_t'(reg2hw.status_503.q);
  assign rcache_line[1][247].status_reg.qe    = reg2hw.status_503.qe;
  assign rcache_line[1][247].status_reg.re    = reg2hw.status_503.re;


  assign rcache_line[1][248].tag_reg.tag      = reg2hw.tag_504.q;
  assign rcache_line[1][248].tag_reg.qe       = reg2hw.tag_504.qe;
  assign rcache_line[1][248].tag_reg.re       = reg2hw.tag_504.re;
  assign rcache_line[1][248].status_reg.status = reg2hw.status_504.q;//status_reg_t'(reg2hw.status_504.q);
  assign rcache_line[1][248].status_reg.qe    = reg2hw.status_504.qe;
  assign rcache_line[1][248].status_reg.re    = reg2hw.status_504.re;


  assign rcache_line[1][249].tag_reg.tag      = reg2hw.tag_505.q;
  assign rcache_line[1][249].tag_reg.qe       = reg2hw.tag_505.qe;
  assign rcache_line[1][249].tag_reg.re       = reg2hw.tag_505.re;
  assign rcache_line[1][249].status_reg.status = reg2hw.status_505.q;//status_reg_t'(reg2hw.status_505.q);
  assign rcache_line[1][249].status_reg.qe    = reg2hw.status_505.qe;
  assign rcache_line[1][249].status_reg.re    = reg2hw.status_505.re;


  assign rcache_line[1][250].tag_reg.tag      = reg2hw.tag_506.q;
  assign rcache_line[1][250].tag_reg.qe       = reg2hw.tag_506.qe;
  assign rcache_line[1][250].tag_reg.re       = reg2hw.tag_506.re;
  assign rcache_line[1][250].status_reg.status = reg2hw.status_506.q;//status_reg_t'(reg2hw.status_506.q);
  assign rcache_line[1][250].status_reg.qe    = reg2hw.status_506.qe;
  assign rcache_line[1][250].status_reg.re    = reg2hw.status_506.re;


  assign rcache_line[1][251].tag_reg.tag      = reg2hw.tag_507.q;
  assign rcache_line[1][251].tag_reg.qe       = reg2hw.tag_507.qe;
  assign rcache_line[1][251].tag_reg.re       = reg2hw.tag_507.re;
  assign rcache_line[1][251].status_reg.status = reg2hw.status_507.q;//status_reg_t'(reg2hw.status_507.q);
  assign rcache_line[1][251].status_reg.qe    = reg2hw.status_507.qe;
  assign rcache_line[1][251].status_reg.re    = reg2hw.status_507.re;


  assign rcache_line[1][252].tag_reg.tag      = reg2hw.tag_508.q;
  assign rcache_line[1][252].tag_reg.qe       = reg2hw.tag_508.qe;
  assign rcache_line[1][252].tag_reg.re       = reg2hw.tag_508.re;
  assign rcache_line[1][252].status_reg.status = reg2hw.status_508.q;//status_reg_t'(reg2hw.status_508.q);
  assign rcache_line[1][252].status_reg.qe    = reg2hw.status_508.qe;
  assign rcache_line[1][252].status_reg.re    = reg2hw.status_508.re;


  assign rcache_line[1][253].tag_reg.tag      = reg2hw.tag_509.q;
  assign rcache_line[1][253].tag_reg.qe       = reg2hw.tag_509.qe;
  assign rcache_line[1][253].tag_reg.re       = reg2hw.tag_509.re;
  assign rcache_line[1][253].status_reg.status = reg2hw.status_509.q;//status_reg_t'(reg2hw.status_509.q);
  assign rcache_line[1][253].status_reg.qe    = reg2hw.status_509.qe;
  assign rcache_line[1][253].status_reg.re    = reg2hw.status_509.re;


  assign rcache_line[1][254].tag_reg.tag      = reg2hw.tag_510.q;
  assign rcache_line[1][254].tag_reg.qe       = reg2hw.tag_510.qe;
  assign rcache_line[1][254].tag_reg.re       = reg2hw.tag_510.re;
  assign rcache_line[1][254].status_reg.status = reg2hw.status_510.q;//status_reg_t'(reg2hw.status_510.q);
  assign rcache_line[1][254].status_reg.qe    = reg2hw.status_510.qe;
  assign rcache_line[1][254].status_reg.re    = reg2hw.status_510.re;


  assign rcache_line[1][255].tag_reg.tag      = reg2hw.tag_511.q;
  assign rcache_line[1][255].tag_reg.qe       = reg2hw.tag_511.qe;
  assign rcache_line[1][255].tag_reg.re       = reg2hw.tag_511.re;
  assign rcache_line[1][255].status_reg.status = reg2hw.status_511.q;//status_reg_t'(reg2hw.status_511.q);
  assign rcache_line[1][255].status_reg.qe    = reg2hw.status_511.qe;
  assign rcache_line[1][255].status_reg.re    = reg2hw.status_511.re;


  assign rcache_line[2][0].tag_reg.tag      = reg2hw.tag_512.q;
  assign rcache_line[2][0].tag_reg.qe       = reg2hw.tag_512.qe;
  assign rcache_line[2][0].tag_reg.re       = reg2hw.tag_512.re;
  assign rcache_line[2][0].status_reg.status = reg2hw.status_512.q;//status_reg_t'(reg2hw.status_512.q);
  assign rcache_line[2][0].status_reg.qe    = reg2hw.status_512.qe;
  assign rcache_line[2][0].status_reg.re    = reg2hw.status_512.re;


  assign rcache_line[2][1].tag_reg.tag      = reg2hw.tag_513.q;
  assign rcache_line[2][1].tag_reg.qe       = reg2hw.tag_513.qe;
  assign rcache_line[2][1].tag_reg.re       = reg2hw.tag_513.re;
  assign rcache_line[2][1].status_reg.status = reg2hw.status_513.q;//status_reg_t'(reg2hw.status_513.q);
  assign rcache_line[2][1].status_reg.qe    = reg2hw.status_513.qe;
  assign rcache_line[2][1].status_reg.re    = reg2hw.status_513.re;


  assign rcache_line[2][2].tag_reg.tag      = reg2hw.tag_514.q;
  assign rcache_line[2][2].tag_reg.qe       = reg2hw.tag_514.qe;
  assign rcache_line[2][2].tag_reg.re       = reg2hw.tag_514.re;
  assign rcache_line[2][2].status_reg.status = reg2hw.status_514.q;//status_reg_t'(reg2hw.status_514.q);
  assign rcache_line[2][2].status_reg.qe    = reg2hw.status_514.qe;
  assign rcache_line[2][2].status_reg.re    = reg2hw.status_514.re;


  assign rcache_line[2][3].tag_reg.tag      = reg2hw.tag_515.q;
  assign rcache_line[2][3].tag_reg.qe       = reg2hw.tag_515.qe;
  assign rcache_line[2][3].tag_reg.re       = reg2hw.tag_515.re;
  assign rcache_line[2][3].status_reg.status = reg2hw.status_515.q;//status_reg_t'(reg2hw.status_515.q);
  assign rcache_line[2][3].status_reg.qe    = reg2hw.status_515.qe;
  assign rcache_line[2][3].status_reg.re    = reg2hw.status_515.re;


  assign rcache_line[2][4].tag_reg.tag      = reg2hw.tag_516.q;
  assign rcache_line[2][4].tag_reg.qe       = reg2hw.tag_516.qe;
  assign rcache_line[2][4].tag_reg.re       = reg2hw.tag_516.re;
  assign rcache_line[2][4].status_reg.status = reg2hw.status_516.q;//status_reg_t'(reg2hw.status_516.q);
  assign rcache_line[2][4].status_reg.qe    = reg2hw.status_516.qe;
  assign rcache_line[2][4].status_reg.re    = reg2hw.status_516.re;


  assign rcache_line[2][5].tag_reg.tag      = reg2hw.tag_517.q;
  assign rcache_line[2][5].tag_reg.qe       = reg2hw.tag_517.qe;
  assign rcache_line[2][5].tag_reg.re       = reg2hw.tag_517.re;
  assign rcache_line[2][5].status_reg.status = reg2hw.status_517.q;//status_reg_t'(reg2hw.status_517.q);
  assign rcache_line[2][5].status_reg.qe    = reg2hw.status_517.qe;
  assign rcache_line[2][5].status_reg.re    = reg2hw.status_517.re;


  assign rcache_line[2][6].tag_reg.tag      = reg2hw.tag_518.q;
  assign rcache_line[2][6].tag_reg.qe       = reg2hw.tag_518.qe;
  assign rcache_line[2][6].tag_reg.re       = reg2hw.tag_518.re;
  assign rcache_line[2][6].status_reg.status = reg2hw.status_518.q;//status_reg_t'(reg2hw.status_518.q);
  assign rcache_line[2][6].status_reg.qe    = reg2hw.status_518.qe;
  assign rcache_line[2][6].status_reg.re    = reg2hw.status_518.re;


  assign rcache_line[2][7].tag_reg.tag      = reg2hw.tag_519.q;
  assign rcache_line[2][7].tag_reg.qe       = reg2hw.tag_519.qe;
  assign rcache_line[2][7].tag_reg.re       = reg2hw.tag_519.re;
  assign rcache_line[2][7].status_reg.status = reg2hw.status_519.q;//status_reg_t'(reg2hw.status_519.q);
  assign rcache_line[2][7].status_reg.qe    = reg2hw.status_519.qe;
  assign rcache_line[2][7].status_reg.re    = reg2hw.status_519.re;


  assign rcache_line[2][8].tag_reg.tag      = reg2hw.tag_520.q;
  assign rcache_line[2][8].tag_reg.qe       = reg2hw.tag_520.qe;
  assign rcache_line[2][8].tag_reg.re       = reg2hw.tag_520.re;
  assign rcache_line[2][8].status_reg.status = reg2hw.status_520.q;//status_reg_t'(reg2hw.status_520.q);
  assign rcache_line[2][8].status_reg.qe    = reg2hw.status_520.qe;
  assign rcache_line[2][8].status_reg.re    = reg2hw.status_520.re;


  assign rcache_line[2][9].tag_reg.tag      = reg2hw.tag_521.q;
  assign rcache_line[2][9].tag_reg.qe       = reg2hw.tag_521.qe;
  assign rcache_line[2][9].tag_reg.re       = reg2hw.tag_521.re;
  assign rcache_line[2][9].status_reg.status = reg2hw.status_521.q;//status_reg_t'(reg2hw.status_521.q);
  assign rcache_line[2][9].status_reg.qe    = reg2hw.status_521.qe;
  assign rcache_line[2][9].status_reg.re    = reg2hw.status_521.re;


  assign rcache_line[2][10].tag_reg.tag      = reg2hw.tag_522.q;
  assign rcache_line[2][10].tag_reg.qe       = reg2hw.tag_522.qe;
  assign rcache_line[2][10].tag_reg.re       = reg2hw.tag_522.re;
  assign rcache_line[2][10].status_reg.status = reg2hw.status_522.q;//status_reg_t'(reg2hw.status_522.q);
  assign rcache_line[2][10].status_reg.qe    = reg2hw.status_522.qe;
  assign rcache_line[2][10].status_reg.re    = reg2hw.status_522.re;


  assign rcache_line[2][11].tag_reg.tag      = reg2hw.tag_523.q;
  assign rcache_line[2][11].tag_reg.qe       = reg2hw.tag_523.qe;
  assign rcache_line[2][11].tag_reg.re       = reg2hw.tag_523.re;
  assign rcache_line[2][11].status_reg.status = reg2hw.status_523.q;//status_reg_t'(reg2hw.status_523.q);
  assign rcache_line[2][11].status_reg.qe    = reg2hw.status_523.qe;
  assign rcache_line[2][11].status_reg.re    = reg2hw.status_523.re;


  assign rcache_line[2][12].tag_reg.tag      = reg2hw.tag_524.q;
  assign rcache_line[2][12].tag_reg.qe       = reg2hw.tag_524.qe;
  assign rcache_line[2][12].tag_reg.re       = reg2hw.tag_524.re;
  assign rcache_line[2][12].status_reg.status = reg2hw.status_524.q;//status_reg_t'(reg2hw.status_524.q);
  assign rcache_line[2][12].status_reg.qe    = reg2hw.status_524.qe;
  assign rcache_line[2][12].status_reg.re    = reg2hw.status_524.re;


  assign rcache_line[2][13].tag_reg.tag      = reg2hw.tag_525.q;
  assign rcache_line[2][13].tag_reg.qe       = reg2hw.tag_525.qe;
  assign rcache_line[2][13].tag_reg.re       = reg2hw.tag_525.re;
  assign rcache_line[2][13].status_reg.status = reg2hw.status_525.q;//status_reg_t'(reg2hw.status_525.q);
  assign rcache_line[2][13].status_reg.qe    = reg2hw.status_525.qe;
  assign rcache_line[2][13].status_reg.re    = reg2hw.status_525.re;


  assign rcache_line[2][14].tag_reg.tag      = reg2hw.tag_526.q;
  assign rcache_line[2][14].tag_reg.qe       = reg2hw.tag_526.qe;
  assign rcache_line[2][14].tag_reg.re       = reg2hw.tag_526.re;
  assign rcache_line[2][14].status_reg.status = reg2hw.status_526.q;//status_reg_t'(reg2hw.status_526.q);
  assign rcache_line[2][14].status_reg.qe    = reg2hw.status_526.qe;
  assign rcache_line[2][14].status_reg.re    = reg2hw.status_526.re;


  assign rcache_line[2][15].tag_reg.tag      = reg2hw.tag_527.q;
  assign rcache_line[2][15].tag_reg.qe       = reg2hw.tag_527.qe;
  assign rcache_line[2][15].tag_reg.re       = reg2hw.tag_527.re;
  assign rcache_line[2][15].status_reg.status = reg2hw.status_527.q;//status_reg_t'(reg2hw.status_527.q);
  assign rcache_line[2][15].status_reg.qe    = reg2hw.status_527.qe;
  assign rcache_line[2][15].status_reg.re    = reg2hw.status_527.re;


  assign rcache_line[2][16].tag_reg.tag      = reg2hw.tag_528.q;
  assign rcache_line[2][16].tag_reg.qe       = reg2hw.tag_528.qe;
  assign rcache_line[2][16].tag_reg.re       = reg2hw.tag_528.re;
  assign rcache_line[2][16].status_reg.status = reg2hw.status_528.q;//status_reg_t'(reg2hw.status_528.q);
  assign rcache_line[2][16].status_reg.qe    = reg2hw.status_528.qe;
  assign rcache_line[2][16].status_reg.re    = reg2hw.status_528.re;


  assign rcache_line[2][17].tag_reg.tag      = reg2hw.tag_529.q;
  assign rcache_line[2][17].tag_reg.qe       = reg2hw.tag_529.qe;
  assign rcache_line[2][17].tag_reg.re       = reg2hw.tag_529.re;
  assign rcache_line[2][17].status_reg.status = reg2hw.status_529.q;//status_reg_t'(reg2hw.status_529.q);
  assign rcache_line[2][17].status_reg.qe    = reg2hw.status_529.qe;
  assign rcache_line[2][17].status_reg.re    = reg2hw.status_529.re;


  assign rcache_line[2][18].tag_reg.tag      = reg2hw.tag_530.q;
  assign rcache_line[2][18].tag_reg.qe       = reg2hw.tag_530.qe;
  assign rcache_line[2][18].tag_reg.re       = reg2hw.tag_530.re;
  assign rcache_line[2][18].status_reg.status = reg2hw.status_530.q;//status_reg_t'(reg2hw.status_530.q);
  assign rcache_line[2][18].status_reg.qe    = reg2hw.status_530.qe;
  assign rcache_line[2][18].status_reg.re    = reg2hw.status_530.re;


  assign rcache_line[2][19].tag_reg.tag      = reg2hw.tag_531.q;
  assign rcache_line[2][19].tag_reg.qe       = reg2hw.tag_531.qe;
  assign rcache_line[2][19].tag_reg.re       = reg2hw.tag_531.re;
  assign rcache_line[2][19].status_reg.status = reg2hw.status_531.q;//status_reg_t'(reg2hw.status_531.q);
  assign rcache_line[2][19].status_reg.qe    = reg2hw.status_531.qe;
  assign rcache_line[2][19].status_reg.re    = reg2hw.status_531.re;


  assign rcache_line[2][20].tag_reg.tag      = reg2hw.tag_532.q;
  assign rcache_line[2][20].tag_reg.qe       = reg2hw.tag_532.qe;
  assign rcache_line[2][20].tag_reg.re       = reg2hw.tag_532.re;
  assign rcache_line[2][20].status_reg.status = reg2hw.status_532.q;//status_reg_t'(reg2hw.status_532.q);
  assign rcache_line[2][20].status_reg.qe    = reg2hw.status_532.qe;
  assign rcache_line[2][20].status_reg.re    = reg2hw.status_532.re;


  assign rcache_line[2][21].tag_reg.tag      = reg2hw.tag_533.q;
  assign rcache_line[2][21].tag_reg.qe       = reg2hw.tag_533.qe;
  assign rcache_line[2][21].tag_reg.re       = reg2hw.tag_533.re;
  assign rcache_line[2][21].status_reg.status = reg2hw.status_533.q;//status_reg_t'(reg2hw.status_533.q);
  assign rcache_line[2][21].status_reg.qe    = reg2hw.status_533.qe;
  assign rcache_line[2][21].status_reg.re    = reg2hw.status_533.re;


  assign rcache_line[2][22].tag_reg.tag      = reg2hw.tag_534.q;
  assign rcache_line[2][22].tag_reg.qe       = reg2hw.tag_534.qe;
  assign rcache_line[2][22].tag_reg.re       = reg2hw.tag_534.re;
  assign rcache_line[2][22].status_reg.status = reg2hw.status_534.q;//status_reg_t'(reg2hw.status_534.q);
  assign rcache_line[2][22].status_reg.qe    = reg2hw.status_534.qe;
  assign rcache_line[2][22].status_reg.re    = reg2hw.status_534.re;


  assign rcache_line[2][23].tag_reg.tag      = reg2hw.tag_535.q;
  assign rcache_line[2][23].tag_reg.qe       = reg2hw.tag_535.qe;
  assign rcache_line[2][23].tag_reg.re       = reg2hw.tag_535.re;
  assign rcache_line[2][23].status_reg.status = reg2hw.status_535.q;//status_reg_t'(reg2hw.status_535.q);
  assign rcache_line[2][23].status_reg.qe    = reg2hw.status_535.qe;
  assign rcache_line[2][23].status_reg.re    = reg2hw.status_535.re;


  assign rcache_line[2][24].tag_reg.tag      = reg2hw.tag_536.q;
  assign rcache_line[2][24].tag_reg.qe       = reg2hw.tag_536.qe;
  assign rcache_line[2][24].tag_reg.re       = reg2hw.tag_536.re;
  assign rcache_line[2][24].status_reg.status = reg2hw.status_536.q;//status_reg_t'(reg2hw.status_536.q);
  assign rcache_line[2][24].status_reg.qe    = reg2hw.status_536.qe;
  assign rcache_line[2][24].status_reg.re    = reg2hw.status_536.re;


  assign rcache_line[2][25].tag_reg.tag      = reg2hw.tag_537.q;
  assign rcache_line[2][25].tag_reg.qe       = reg2hw.tag_537.qe;
  assign rcache_line[2][25].tag_reg.re       = reg2hw.tag_537.re;
  assign rcache_line[2][25].status_reg.status = reg2hw.status_537.q;//status_reg_t'(reg2hw.status_537.q);
  assign rcache_line[2][25].status_reg.qe    = reg2hw.status_537.qe;
  assign rcache_line[2][25].status_reg.re    = reg2hw.status_537.re;


  assign rcache_line[2][26].tag_reg.tag      = reg2hw.tag_538.q;
  assign rcache_line[2][26].tag_reg.qe       = reg2hw.tag_538.qe;
  assign rcache_line[2][26].tag_reg.re       = reg2hw.tag_538.re;
  assign rcache_line[2][26].status_reg.status = reg2hw.status_538.q;//status_reg_t'(reg2hw.status_538.q);
  assign rcache_line[2][26].status_reg.qe    = reg2hw.status_538.qe;
  assign rcache_line[2][26].status_reg.re    = reg2hw.status_538.re;


  assign rcache_line[2][27].tag_reg.tag      = reg2hw.tag_539.q;
  assign rcache_line[2][27].tag_reg.qe       = reg2hw.tag_539.qe;
  assign rcache_line[2][27].tag_reg.re       = reg2hw.tag_539.re;
  assign rcache_line[2][27].status_reg.status = reg2hw.status_539.q;//status_reg_t'(reg2hw.status_539.q);
  assign rcache_line[2][27].status_reg.qe    = reg2hw.status_539.qe;
  assign rcache_line[2][27].status_reg.re    = reg2hw.status_539.re;


  assign rcache_line[2][28].tag_reg.tag      = reg2hw.tag_540.q;
  assign rcache_line[2][28].tag_reg.qe       = reg2hw.tag_540.qe;
  assign rcache_line[2][28].tag_reg.re       = reg2hw.tag_540.re;
  assign rcache_line[2][28].status_reg.status = reg2hw.status_540.q;//status_reg_t'(reg2hw.status_540.q);
  assign rcache_line[2][28].status_reg.qe    = reg2hw.status_540.qe;
  assign rcache_line[2][28].status_reg.re    = reg2hw.status_540.re;


  assign rcache_line[2][29].tag_reg.tag      = reg2hw.tag_541.q;
  assign rcache_line[2][29].tag_reg.qe       = reg2hw.tag_541.qe;
  assign rcache_line[2][29].tag_reg.re       = reg2hw.tag_541.re;
  assign rcache_line[2][29].status_reg.status = reg2hw.status_541.q;//status_reg_t'(reg2hw.status_541.q);
  assign rcache_line[2][29].status_reg.qe    = reg2hw.status_541.qe;
  assign rcache_line[2][29].status_reg.re    = reg2hw.status_541.re;


  assign rcache_line[2][30].tag_reg.tag      = reg2hw.tag_542.q;
  assign rcache_line[2][30].tag_reg.qe       = reg2hw.tag_542.qe;
  assign rcache_line[2][30].tag_reg.re       = reg2hw.tag_542.re;
  assign rcache_line[2][30].status_reg.status = reg2hw.status_542.q;//status_reg_t'(reg2hw.status_542.q);
  assign rcache_line[2][30].status_reg.qe    = reg2hw.status_542.qe;
  assign rcache_line[2][30].status_reg.re    = reg2hw.status_542.re;


  assign rcache_line[2][31].tag_reg.tag      = reg2hw.tag_543.q;
  assign rcache_line[2][31].tag_reg.qe       = reg2hw.tag_543.qe;
  assign rcache_line[2][31].tag_reg.re       = reg2hw.tag_543.re;
  assign rcache_line[2][31].status_reg.status = reg2hw.status_543.q;//status_reg_t'(reg2hw.status_543.q);
  assign rcache_line[2][31].status_reg.qe    = reg2hw.status_543.qe;
  assign rcache_line[2][31].status_reg.re    = reg2hw.status_543.re;


  assign rcache_line[2][32].tag_reg.tag      = reg2hw.tag_544.q;
  assign rcache_line[2][32].tag_reg.qe       = reg2hw.tag_544.qe;
  assign rcache_line[2][32].tag_reg.re       = reg2hw.tag_544.re;
  assign rcache_line[2][32].status_reg.status = reg2hw.status_544.q;//status_reg_t'(reg2hw.status_544.q);
  assign rcache_line[2][32].status_reg.qe    = reg2hw.status_544.qe;
  assign rcache_line[2][32].status_reg.re    = reg2hw.status_544.re;


  assign rcache_line[2][33].tag_reg.tag      = reg2hw.tag_545.q;
  assign rcache_line[2][33].tag_reg.qe       = reg2hw.tag_545.qe;
  assign rcache_line[2][33].tag_reg.re       = reg2hw.tag_545.re;
  assign rcache_line[2][33].status_reg.status = reg2hw.status_545.q;//status_reg_t'(reg2hw.status_545.q);
  assign rcache_line[2][33].status_reg.qe    = reg2hw.status_545.qe;
  assign rcache_line[2][33].status_reg.re    = reg2hw.status_545.re;


  assign rcache_line[2][34].tag_reg.tag      = reg2hw.tag_546.q;
  assign rcache_line[2][34].tag_reg.qe       = reg2hw.tag_546.qe;
  assign rcache_line[2][34].tag_reg.re       = reg2hw.tag_546.re;
  assign rcache_line[2][34].status_reg.status = reg2hw.status_546.q;//status_reg_t'(reg2hw.status_546.q);
  assign rcache_line[2][34].status_reg.qe    = reg2hw.status_546.qe;
  assign rcache_line[2][34].status_reg.re    = reg2hw.status_546.re;


  assign rcache_line[2][35].tag_reg.tag      = reg2hw.tag_547.q;
  assign rcache_line[2][35].tag_reg.qe       = reg2hw.tag_547.qe;
  assign rcache_line[2][35].tag_reg.re       = reg2hw.tag_547.re;
  assign rcache_line[2][35].status_reg.status = reg2hw.status_547.q;//status_reg_t'(reg2hw.status_547.q);
  assign rcache_line[2][35].status_reg.qe    = reg2hw.status_547.qe;
  assign rcache_line[2][35].status_reg.re    = reg2hw.status_547.re;


  assign rcache_line[2][36].tag_reg.tag      = reg2hw.tag_548.q;
  assign rcache_line[2][36].tag_reg.qe       = reg2hw.tag_548.qe;
  assign rcache_line[2][36].tag_reg.re       = reg2hw.tag_548.re;
  assign rcache_line[2][36].status_reg.status = reg2hw.status_548.q;//status_reg_t'(reg2hw.status_548.q);
  assign rcache_line[2][36].status_reg.qe    = reg2hw.status_548.qe;
  assign rcache_line[2][36].status_reg.re    = reg2hw.status_548.re;


  assign rcache_line[2][37].tag_reg.tag      = reg2hw.tag_549.q;
  assign rcache_line[2][37].tag_reg.qe       = reg2hw.tag_549.qe;
  assign rcache_line[2][37].tag_reg.re       = reg2hw.tag_549.re;
  assign rcache_line[2][37].status_reg.status = reg2hw.status_549.q;//status_reg_t'(reg2hw.status_549.q);
  assign rcache_line[2][37].status_reg.qe    = reg2hw.status_549.qe;
  assign rcache_line[2][37].status_reg.re    = reg2hw.status_549.re;


  assign rcache_line[2][38].tag_reg.tag      = reg2hw.tag_550.q;
  assign rcache_line[2][38].tag_reg.qe       = reg2hw.tag_550.qe;
  assign rcache_line[2][38].tag_reg.re       = reg2hw.tag_550.re;
  assign rcache_line[2][38].status_reg.status = reg2hw.status_550.q;//status_reg_t'(reg2hw.status_550.q);
  assign rcache_line[2][38].status_reg.qe    = reg2hw.status_550.qe;
  assign rcache_line[2][38].status_reg.re    = reg2hw.status_550.re;


  assign rcache_line[2][39].tag_reg.tag      = reg2hw.tag_551.q;
  assign rcache_line[2][39].tag_reg.qe       = reg2hw.tag_551.qe;
  assign rcache_line[2][39].tag_reg.re       = reg2hw.tag_551.re;
  assign rcache_line[2][39].status_reg.status = reg2hw.status_551.q;//status_reg_t'(reg2hw.status_551.q);
  assign rcache_line[2][39].status_reg.qe    = reg2hw.status_551.qe;
  assign rcache_line[2][39].status_reg.re    = reg2hw.status_551.re;


  assign rcache_line[2][40].tag_reg.tag      = reg2hw.tag_552.q;
  assign rcache_line[2][40].tag_reg.qe       = reg2hw.tag_552.qe;
  assign rcache_line[2][40].tag_reg.re       = reg2hw.tag_552.re;
  assign rcache_line[2][40].status_reg.status = reg2hw.status_552.q;//status_reg_t'(reg2hw.status_552.q);
  assign rcache_line[2][40].status_reg.qe    = reg2hw.status_552.qe;
  assign rcache_line[2][40].status_reg.re    = reg2hw.status_552.re;


  assign rcache_line[2][41].tag_reg.tag      = reg2hw.tag_553.q;
  assign rcache_line[2][41].tag_reg.qe       = reg2hw.tag_553.qe;
  assign rcache_line[2][41].tag_reg.re       = reg2hw.tag_553.re;
  assign rcache_line[2][41].status_reg.status = reg2hw.status_553.q;//status_reg_t'(reg2hw.status_553.q);
  assign rcache_line[2][41].status_reg.qe    = reg2hw.status_553.qe;
  assign rcache_line[2][41].status_reg.re    = reg2hw.status_553.re;


  assign rcache_line[2][42].tag_reg.tag      = reg2hw.tag_554.q;
  assign rcache_line[2][42].tag_reg.qe       = reg2hw.tag_554.qe;
  assign rcache_line[2][42].tag_reg.re       = reg2hw.tag_554.re;
  assign rcache_line[2][42].status_reg.status = reg2hw.status_554.q;//status_reg_t'(reg2hw.status_554.q);
  assign rcache_line[2][42].status_reg.qe    = reg2hw.status_554.qe;
  assign rcache_line[2][42].status_reg.re    = reg2hw.status_554.re;


  assign rcache_line[2][43].tag_reg.tag      = reg2hw.tag_555.q;
  assign rcache_line[2][43].tag_reg.qe       = reg2hw.tag_555.qe;
  assign rcache_line[2][43].tag_reg.re       = reg2hw.tag_555.re;
  assign rcache_line[2][43].status_reg.status = reg2hw.status_555.q;//status_reg_t'(reg2hw.status_555.q);
  assign rcache_line[2][43].status_reg.qe    = reg2hw.status_555.qe;
  assign rcache_line[2][43].status_reg.re    = reg2hw.status_555.re;


  assign rcache_line[2][44].tag_reg.tag      = reg2hw.tag_556.q;
  assign rcache_line[2][44].tag_reg.qe       = reg2hw.tag_556.qe;
  assign rcache_line[2][44].tag_reg.re       = reg2hw.tag_556.re;
  assign rcache_line[2][44].status_reg.status = reg2hw.status_556.q;//status_reg_t'(reg2hw.status_556.q);
  assign rcache_line[2][44].status_reg.qe    = reg2hw.status_556.qe;
  assign rcache_line[2][44].status_reg.re    = reg2hw.status_556.re;


  assign rcache_line[2][45].tag_reg.tag      = reg2hw.tag_557.q;
  assign rcache_line[2][45].tag_reg.qe       = reg2hw.tag_557.qe;
  assign rcache_line[2][45].tag_reg.re       = reg2hw.tag_557.re;
  assign rcache_line[2][45].status_reg.status = reg2hw.status_557.q;//status_reg_t'(reg2hw.status_557.q);
  assign rcache_line[2][45].status_reg.qe    = reg2hw.status_557.qe;
  assign rcache_line[2][45].status_reg.re    = reg2hw.status_557.re;


  assign rcache_line[2][46].tag_reg.tag      = reg2hw.tag_558.q;
  assign rcache_line[2][46].tag_reg.qe       = reg2hw.tag_558.qe;
  assign rcache_line[2][46].tag_reg.re       = reg2hw.tag_558.re;
  assign rcache_line[2][46].status_reg.status = reg2hw.status_558.q;//status_reg_t'(reg2hw.status_558.q);
  assign rcache_line[2][46].status_reg.qe    = reg2hw.status_558.qe;
  assign rcache_line[2][46].status_reg.re    = reg2hw.status_558.re;


  assign rcache_line[2][47].tag_reg.tag      = reg2hw.tag_559.q;
  assign rcache_line[2][47].tag_reg.qe       = reg2hw.tag_559.qe;
  assign rcache_line[2][47].tag_reg.re       = reg2hw.tag_559.re;
  assign rcache_line[2][47].status_reg.status = reg2hw.status_559.q;//status_reg_t'(reg2hw.status_559.q);
  assign rcache_line[2][47].status_reg.qe    = reg2hw.status_559.qe;
  assign rcache_line[2][47].status_reg.re    = reg2hw.status_559.re;


  assign rcache_line[2][48].tag_reg.tag      = reg2hw.tag_560.q;
  assign rcache_line[2][48].tag_reg.qe       = reg2hw.tag_560.qe;
  assign rcache_line[2][48].tag_reg.re       = reg2hw.tag_560.re;
  assign rcache_line[2][48].status_reg.status = reg2hw.status_560.q;//status_reg_t'(reg2hw.status_560.q);
  assign rcache_line[2][48].status_reg.qe    = reg2hw.status_560.qe;
  assign rcache_line[2][48].status_reg.re    = reg2hw.status_560.re;


  assign rcache_line[2][49].tag_reg.tag      = reg2hw.tag_561.q;
  assign rcache_line[2][49].tag_reg.qe       = reg2hw.tag_561.qe;
  assign rcache_line[2][49].tag_reg.re       = reg2hw.tag_561.re;
  assign rcache_line[2][49].status_reg.status = reg2hw.status_561.q;//status_reg_t'(reg2hw.status_561.q);
  assign rcache_line[2][49].status_reg.qe    = reg2hw.status_561.qe;
  assign rcache_line[2][49].status_reg.re    = reg2hw.status_561.re;


  assign rcache_line[2][50].tag_reg.tag      = reg2hw.tag_562.q;
  assign rcache_line[2][50].tag_reg.qe       = reg2hw.tag_562.qe;
  assign rcache_line[2][50].tag_reg.re       = reg2hw.tag_562.re;
  assign rcache_line[2][50].status_reg.status = reg2hw.status_562.q;//status_reg_t'(reg2hw.status_562.q);
  assign rcache_line[2][50].status_reg.qe    = reg2hw.status_562.qe;
  assign rcache_line[2][50].status_reg.re    = reg2hw.status_562.re;


  assign rcache_line[2][51].tag_reg.tag      = reg2hw.tag_563.q;
  assign rcache_line[2][51].tag_reg.qe       = reg2hw.tag_563.qe;
  assign rcache_line[2][51].tag_reg.re       = reg2hw.tag_563.re;
  assign rcache_line[2][51].status_reg.status = reg2hw.status_563.q;//status_reg_t'(reg2hw.status_563.q);
  assign rcache_line[2][51].status_reg.qe    = reg2hw.status_563.qe;
  assign rcache_line[2][51].status_reg.re    = reg2hw.status_563.re;


  assign rcache_line[2][52].tag_reg.tag      = reg2hw.tag_564.q;
  assign rcache_line[2][52].tag_reg.qe       = reg2hw.tag_564.qe;
  assign rcache_line[2][52].tag_reg.re       = reg2hw.tag_564.re;
  assign rcache_line[2][52].status_reg.status = reg2hw.status_564.q;//status_reg_t'(reg2hw.status_564.q);
  assign rcache_line[2][52].status_reg.qe    = reg2hw.status_564.qe;
  assign rcache_line[2][52].status_reg.re    = reg2hw.status_564.re;


  assign rcache_line[2][53].tag_reg.tag      = reg2hw.tag_565.q;
  assign rcache_line[2][53].tag_reg.qe       = reg2hw.tag_565.qe;
  assign rcache_line[2][53].tag_reg.re       = reg2hw.tag_565.re;
  assign rcache_line[2][53].status_reg.status = reg2hw.status_565.q;//status_reg_t'(reg2hw.status_565.q);
  assign rcache_line[2][53].status_reg.qe    = reg2hw.status_565.qe;
  assign rcache_line[2][53].status_reg.re    = reg2hw.status_565.re;


  assign rcache_line[2][54].tag_reg.tag      = reg2hw.tag_566.q;
  assign rcache_line[2][54].tag_reg.qe       = reg2hw.tag_566.qe;
  assign rcache_line[2][54].tag_reg.re       = reg2hw.tag_566.re;
  assign rcache_line[2][54].status_reg.status = reg2hw.status_566.q;//status_reg_t'(reg2hw.status_566.q);
  assign rcache_line[2][54].status_reg.qe    = reg2hw.status_566.qe;
  assign rcache_line[2][54].status_reg.re    = reg2hw.status_566.re;


  assign rcache_line[2][55].tag_reg.tag      = reg2hw.tag_567.q;
  assign rcache_line[2][55].tag_reg.qe       = reg2hw.tag_567.qe;
  assign rcache_line[2][55].tag_reg.re       = reg2hw.tag_567.re;
  assign rcache_line[2][55].status_reg.status = reg2hw.status_567.q;//status_reg_t'(reg2hw.status_567.q);
  assign rcache_line[2][55].status_reg.qe    = reg2hw.status_567.qe;
  assign rcache_line[2][55].status_reg.re    = reg2hw.status_567.re;


  assign rcache_line[2][56].tag_reg.tag      = reg2hw.tag_568.q;
  assign rcache_line[2][56].tag_reg.qe       = reg2hw.tag_568.qe;
  assign rcache_line[2][56].tag_reg.re       = reg2hw.tag_568.re;
  assign rcache_line[2][56].status_reg.status = reg2hw.status_568.q;//status_reg_t'(reg2hw.status_568.q);
  assign rcache_line[2][56].status_reg.qe    = reg2hw.status_568.qe;
  assign rcache_line[2][56].status_reg.re    = reg2hw.status_568.re;


  assign rcache_line[2][57].tag_reg.tag      = reg2hw.tag_569.q;
  assign rcache_line[2][57].tag_reg.qe       = reg2hw.tag_569.qe;
  assign rcache_line[2][57].tag_reg.re       = reg2hw.tag_569.re;
  assign rcache_line[2][57].status_reg.status = reg2hw.status_569.q;//status_reg_t'(reg2hw.status_569.q);
  assign rcache_line[2][57].status_reg.qe    = reg2hw.status_569.qe;
  assign rcache_line[2][57].status_reg.re    = reg2hw.status_569.re;


  assign rcache_line[2][58].tag_reg.tag      = reg2hw.tag_570.q;
  assign rcache_line[2][58].tag_reg.qe       = reg2hw.tag_570.qe;
  assign rcache_line[2][58].tag_reg.re       = reg2hw.tag_570.re;
  assign rcache_line[2][58].status_reg.status = reg2hw.status_570.q;//status_reg_t'(reg2hw.status_570.q);
  assign rcache_line[2][58].status_reg.qe    = reg2hw.status_570.qe;
  assign rcache_line[2][58].status_reg.re    = reg2hw.status_570.re;


  assign rcache_line[2][59].tag_reg.tag      = reg2hw.tag_571.q;
  assign rcache_line[2][59].tag_reg.qe       = reg2hw.tag_571.qe;
  assign rcache_line[2][59].tag_reg.re       = reg2hw.tag_571.re;
  assign rcache_line[2][59].status_reg.status = reg2hw.status_571.q;//status_reg_t'(reg2hw.status_571.q);
  assign rcache_line[2][59].status_reg.qe    = reg2hw.status_571.qe;
  assign rcache_line[2][59].status_reg.re    = reg2hw.status_571.re;


  assign rcache_line[2][60].tag_reg.tag      = reg2hw.tag_572.q;
  assign rcache_line[2][60].tag_reg.qe       = reg2hw.tag_572.qe;
  assign rcache_line[2][60].tag_reg.re       = reg2hw.tag_572.re;
  assign rcache_line[2][60].status_reg.status = reg2hw.status_572.q;//status_reg_t'(reg2hw.status_572.q);
  assign rcache_line[2][60].status_reg.qe    = reg2hw.status_572.qe;
  assign rcache_line[2][60].status_reg.re    = reg2hw.status_572.re;


  assign rcache_line[2][61].tag_reg.tag      = reg2hw.tag_573.q;
  assign rcache_line[2][61].tag_reg.qe       = reg2hw.tag_573.qe;
  assign rcache_line[2][61].tag_reg.re       = reg2hw.tag_573.re;
  assign rcache_line[2][61].status_reg.status = reg2hw.status_573.q;//status_reg_t'(reg2hw.status_573.q);
  assign rcache_line[2][61].status_reg.qe    = reg2hw.status_573.qe;
  assign rcache_line[2][61].status_reg.re    = reg2hw.status_573.re;


  assign rcache_line[2][62].tag_reg.tag      = reg2hw.tag_574.q;
  assign rcache_line[2][62].tag_reg.qe       = reg2hw.tag_574.qe;
  assign rcache_line[2][62].tag_reg.re       = reg2hw.tag_574.re;
  assign rcache_line[2][62].status_reg.status = reg2hw.status_574.q;//status_reg_t'(reg2hw.status_574.q);
  assign rcache_line[2][62].status_reg.qe    = reg2hw.status_574.qe;
  assign rcache_line[2][62].status_reg.re    = reg2hw.status_574.re;


  assign rcache_line[2][63].tag_reg.tag      = reg2hw.tag_575.q;
  assign rcache_line[2][63].tag_reg.qe       = reg2hw.tag_575.qe;
  assign rcache_line[2][63].tag_reg.re       = reg2hw.tag_575.re;
  assign rcache_line[2][63].status_reg.status = reg2hw.status_575.q;//status_reg_t'(reg2hw.status_575.q);
  assign rcache_line[2][63].status_reg.qe    = reg2hw.status_575.qe;
  assign rcache_line[2][63].status_reg.re    = reg2hw.status_575.re;


  assign rcache_line[2][64].tag_reg.tag      = reg2hw.tag_576.q;
  assign rcache_line[2][64].tag_reg.qe       = reg2hw.tag_576.qe;
  assign rcache_line[2][64].tag_reg.re       = reg2hw.tag_576.re;
  assign rcache_line[2][64].status_reg.status = reg2hw.status_576.q;//status_reg_t'(reg2hw.status_576.q);
  assign rcache_line[2][64].status_reg.qe    = reg2hw.status_576.qe;
  assign rcache_line[2][64].status_reg.re    = reg2hw.status_576.re;


  assign rcache_line[2][65].tag_reg.tag      = reg2hw.tag_577.q;
  assign rcache_line[2][65].tag_reg.qe       = reg2hw.tag_577.qe;
  assign rcache_line[2][65].tag_reg.re       = reg2hw.tag_577.re;
  assign rcache_line[2][65].status_reg.status = reg2hw.status_577.q;//status_reg_t'(reg2hw.status_577.q);
  assign rcache_line[2][65].status_reg.qe    = reg2hw.status_577.qe;
  assign rcache_line[2][65].status_reg.re    = reg2hw.status_577.re;


  assign rcache_line[2][66].tag_reg.tag      = reg2hw.tag_578.q;
  assign rcache_line[2][66].tag_reg.qe       = reg2hw.tag_578.qe;
  assign rcache_line[2][66].tag_reg.re       = reg2hw.tag_578.re;
  assign rcache_line[2][66].status_reg.status = reg2hw.status_578.q;//status_reg_t'(reg2hw.status_578.q);
  assign rcache_line[2][66].status_reg.qe    = reg2hw.status_578.qe;
  assign rcache_line[2][66].status_reg.re    = reg2hw.status_578.re;


  assign rcache_line[2][67].tag_reg.tag      = reg2hw.tag_579.q;
  assign rcache_line[2][67].tag_reg.qe       = reg2hw.tag_579.qe;
  assign rcache_line[2][67].tag_reg.re       = reg2hw.tag_579.re;
  assign rcache_line[2][67].status_reg.status = reg2hw.status_579.q;//status_reg_t'(reg2hw.status_579.q);
  assign rcache_line[2][67].status_reg.qe    = reg2hw.status_579.qe;
  assign rcache_line[2][67].status_reg.re    = reg2hw.status_579.re;


  assign rcache_line[2][68].tag_reg.tag      = reg2hw.tag_580.q;
  assign rcache_line[2][68].tag_reg.qe       = reg2hw.tag_580.qe;
  assign rcache_line[2][68].tag_reg.re       = reg2hw.tag_580.re;
  assign rcache_line[2][68].status_reg.status = reg2hw.status_580.q;//status_reg_t'(reg2hw.status_580.q);
  assign rcache_line[2][68].status_reg.qe    = reg2hw.status_580.qe;
  assign rcache_line[2][68].status_reg.re    = reg2hw.status_580.re;


  assign rcache_line[2][69].tag_reg.tag      = reg2hw.tag_581.q;
  assign rcache_line[2][69].tag_reg.qe       = reg2hw.tag_581.qe;
  assign rcache_line[2][69].tag_reg.re       = reg2hw.tag_581.re;
  assign rcache_line[2][69].status_reg.status = reg2hw.status_581.q;//status_reg_t'(reg2hw.status_581.q);
  assign rcache_line[2][69].status_reg.qe    = reg2hw.status_581.qe;
  assign rcache_line[2][69].status_reg.re    = reg2hw.status_581.re;


  assign rcache_line[2][70].tag_reg.tag      = reg2hw.tag_582.q;
  assign rcache_line[2][70].tag_reg.qe       = reg2hw.tag_582.qe;
  assign rcache_line[2][70].tag_reg.re       = reg2hw.tag_582.re;
  assign rcache_line[2][70].status_reg.status = reg2hw.status_582.q;//status_reg_t'(reg2hw.status_582.q);
  assign rcache_line[2][70].status_reg.qe    = reg2hw.status_582.qe;
  assign rcache_line[2][70].status_reg.re    = reg2hw.status_582.re;


  assign rcache_line[2][71].tag_reg.tag      = reg2hw.tag_583.q;
  assign rcache_line[2][71].tag_reg.qe       = reg2hw.tag_583.qe;
  assign rcache_line[2][71].tag_reg.re       = reg2hw.tag_583.re;
  assign rcache_line[2][71].status_reg.status = reg2hw.status_583.q;//status_reg_t'(reg2hw.status_583.q);
  assign rcache_line[2][71].status_reg.qe    = reg2hw.status_583.qe;
  assign rcache_line[2][71].status_reg.re    = reg2hw.status_583.re;


  assign rcache_line[2][72].tag_reg.tag      = reg2hw.tag_584.q;
  assign rcache_line[2][72].tag_reg.qe       = reg2hw.tag_584.qe;
  assign rcache_line[2][72].tag_reg.re       = reg2hw.tag_584.re;
  assign rcache_line[2][72].status_reg.status = reg2hw.status_584.q;//status_reg_t'(reg2hw.status_584.q);
  assign rcache_line[2][72].status_reg.qe    = reg2hw.status_584.qe;
  assign rcache_line[2][72].status_reg.re    = reg2hw.status_584.re;


  assign rcache_line[2][73].tag_reg.tag      = reg2hw.tag_585.q;
  assign rcache_line[2][73].tag_reg.qe       = reg2hw.tag_585.qe;
  assign rcache_line[2][73].tag_reg.re       = reg2hw.tag_585.re;
  assign rcache_line[2][73].status_reg.status = reg2hw.status_585.q;//status_reg_t'(reg2hw.status_585.q);
  assign rcache_line[2][73].status_reg.qe    = reg2hw.status_585.qe;
  assign rcache_line[2][73].status_reg.re    = reg2hw.status_585.re;


  assign rcache_line[2][74].tag_reg.tag      = reg2hw.tag_586.q;
  assign rcache_line[2][74].tag_reg.qe       = reg2hw.tag_586.qe;
  assign rcache_line[2][74].tag_reg.re       = reg2hw.tag_586.re;
  assign rcache_line[2][74].status_reg.status = reg2hw.status_586.q;//status_reg_t'(reg2hw.status_586.q);
  assign rcache_line[2][74].status_reg.qe    = reg2hw.status_586.qe;
  assign rcache_line[2][74].status_reg.re    = reg2hw.status_586.re;


  assign rcache_line[2][75].tag_reg.tag      = reg2hw.tag_587.q;
  assign rcache_line[2][75].tag_reg.qe       = reg2hw.tag_587.qe;
  assign rcache_line[2][75].tag_reg.re       = reg2hw.tag_587.re;
  assign rcache_line[2][75].status_reg.status = reg2hw.status_587.q;//status_reg_t'(reg2hw.status_587.q);
  assign rcache_line[2][75].status_reg.qe    = reg2hw.status_587.qe;
  assign rcache_line[2][75].status_reg.re    = reg2hw.status_587.re;


  assign rcache_line[2][76].tag_reg.tag      = reg2hw.tag_588.q;
  assign rcache_line[2][76].tag_reg.qe       = reg2hw.tag_588.qe;
  assign rcache_line[2][76].tag_reg.re       = reg2hw.tag_588.re;
  assign rcache_line[2][76].status_reg.status = reg2hw.status_588.q;//status_reg_t'(reg2hw.status_588.q);
  assign rcache_line[2][76].status_reg.qe    = reg2hw.status_588.qe;
  assign rcache_line[2][76].status_reg.re    = reg2hw.status_588.re;


  assign rcache_line[2][77].tag_reg.tag      = reg2hw.tag_589.q;
  assign rcache_line[2][77].tag_reg.qe       = reg2hw.tag_589.qe;
  assign rcache_line[2][77].tag_reg.re       = reg2hw.tag_589.re;
  assign rcache_line[2][77].status_reg.status = reg2hw.status_589.q;//status_reg_t'(reg2hw.status_589.q);
  assign rcache_line[2][77].status_reg.qe    = reg2hw.status_589.qe;
  assign rcache_line[2][77].status_reg.re    = reg2hw.status_589.re;


  assign rcache_line[2][78].tag_reg.tag      = reg2hw.tag_590.q;
  assign rcache_line[2][78].tag_reg.qe       = reg2hw.tag_590.qe;
  assign rcache_line[2][78].tag_reg.re       = reg2hw.tag_590.re;
  assign rcache_line[2][78].status_reg.status = reg2hw.status_590.q;//status_reg_t'(reg2hw.status_590.q);
  assign rcache_line[2][78].status_reg.qe    = reg2hw.status_590.qe;
  assign rcache_line[2][78].status_reg.re    = reg2hw.status_590.re;


  assign rcache_line[2][79].tag_reg.tag      = reg2hw.tag_591.q;
  assign rcache_line[2][79].tag_reg.qe       = reg2hw.tag_591.qe;
  assign rcache_line[2][79].tag_reg.re       = reg2hw.tag_591.re;
  assign rcache_line[2][79].status_reg.status = reg2hw.status_591.q;//status_reg_t'(reg2hw.status_591.q);
  assign rcache_line[2][79].status_reg.qe    = reg2hw.status_591.qe;
  assign rcache_line[2][79].status_reg.re    = reg2hw.status_591.re;


  assign rcache_line[2][80].tag_reg.tag      = reg2hw.tag_592.q;
  assign rcache_line[2][80].tag_reg.qe       = reg2hw.tag_592.qe;
  assign rcache_line[2][80].tag_reg.re       = reg2hw.tag_592.re;
  assign rcache_line[2][80].status_reg.status = reg2hw.status_592.q;//status_reg_t'(reg2hw.status_592.q);
  assign rcache_line[2][80].status_reg.qe    = reg2hw.status_592.qe;
  assign rcache_line[2][80].status_reg.re    = reg2hw.status_592.re;


  assign rcache_line[2][81].tag_reg.tag      = reg2hw.tag_593.q;
  assign rcache_line[2][81].tag_reg.qe       = reg2hw.tag_593.qe;
  assign rcache_line[2][81].tag_reg.re       = reg2hw.tag_593.re;
  assign rcache_line[2][81].status_reg.status = reg2hw.status_593.q;//status_reg_t'(reg2hw.status_593.q);
  assign rcache_line[2][81].status_reg.qe    = reg2hw.status_593.qe;
  assign rcache_line[2][81].status_reg.re    = reg2hw.status_593.re;


  assign rcache_line[2][82].tag_reg.tag      = reg2hw.tag_594.q;
  assign rcache_line[2][82].tag_reg.qe       = reg2hw.tag_594.qe;
  assign rcache_line[2][82].tag_reg.re       = reg2hw.tag_594.re;
  assign rcache_line[2][82].status_reg.status = reg2hw.status_594.q;//status_reg_t'(reg2hw.status_594.q);
  assign rcache_line[2][82].status_reg.qe    = reg2hw.status_594.qe;
  assign rcache_line[2][82].status_reg.re    = reg2hw.status_594.re;


  assign rcache_line[2][83].tag_reg.tag      = reg2hw.tag_595.q;
  assign rcache_line[2][83].tag_reg.qe       = reg2hw.tag_595.qe;
  assign rcache_line[2][83].tag_reg.re       = reg2hw.tag_595.re;
  assign rcache_line[2][83].status_reg.status = reg2hw.status_595.q;//status_reg_t'(reg2hw.status_595.q);
  assign rcache_line[2][83].status_reg.qe    = reg2hw.status_595.qe;
  assign rcache_line[2][83].status_reg.re    = reg2hw.status_595.re;


  assign rcache_line[2][84].tag_reg.tag      = reg2hw.tag_596.q;
  assign rcache_line[2][84].tag_reg.qe       = reg2hw.tag_596.qe;
  assign rcache_line[2][84].tag_reg.re       = reg2hw.tag_596.re;
  assign rcache_line[2][84].status_reg.status = reg2hw.status_596.q;//status_reg_t'(reg2hw.status_596.q);
  assign rcache_line[2][84].status_reg.qe    = reg2hw.status_596.qe;
  assign rcache_line[2][84].status_reg.re    = reg2hw.status_596.re;


  assign rcache_line[2][85].tag_reg.tag      = reg2hw.tag_597.q;
  assign rcache_line[2][85].tag_reg.qe       = reg2hw.tag_597.qe;
  assign rcache_line[2][85].tag_reg.re       = reg2hw.tag_597.re;
  assign rcache_line[2][85].status_reg.status = reg2hw.status_597.q;//status_reg_t'(reg2hw.status_597.q);
  assign rcache_line[2][85].status_reg.qe    = reg2hw.status_597.qe;
  assign rcache_line[2][85].status_reg.re    = reg2hw.status_597.re;


  assign rcache_line[2][86].tag_reg.tag      = reg2hw.tag_598.q;
  assign rcache_line[2][86].tag_reg.qe       = reg2hw.tag_598.qe;
  assign rcache_line[2][86].tag_reg.re       = reg2hw.tag_598.re;
  assign rcache_line[2][86].status_reg.status = reg2hw.status_598.q;//status_reg_t'(reg2hw.status_598.q);
  assign rcache_line[2][86].status_reg.qe    = reg2hw.status_598.qe;
  assign rcache_line[2][86].status_reg.re    = reg2hw.status_598.re;


  assign rcache_line[2][87].tag_reg.tag      = reg2hw.tag_599.q;
  assign rcache_line[2][87].tag_reg.qe       = reg2hw.tag_599.qe;
  assign rcache_line[2][87].tag_reg.re       = reg2hw.tag_599.re;
  assign rcache_line[2][87].status_reg.status = reg2hw.status_599.q;//status_reg_t'(reg2hw.status_599.q);
  assign rcache_line[2][87].status_reg.qe    = reg2hw.status_599.qe;
  assign rcache_line[2][87].status_reg.re    = reg2hw.status_599.re;


  assign rcache_line[2][88].tag_reg.tag      = reg2hw.tag_600.q;
  assign rcache_line[2][88].tag_reg.qe       = reg2hw.tag_600.qe;
  assign rcache_line[2][88].tag_reg.re       = reg2hw.tag_600.re;
  assign rcache_line[2][88].status_reg.status = reg2hw.status_600.q;//status_reg_t'(reg2hw.status_600.q);
  assign rcache_line[2][88].status_reg.qe    = reg2hw.status_600.qe;
  assign rcache_line[2][88].status_reg.re    = reg2hw.status_600.re;


  assign rcache_line[2][89].tag_reg.tag      = reg2hw.tag_601.q;
  assign rcache_line[2][89].tag_reg.qe       = reg2hw.tag_601.qe;
  assign rcache_line[2][89].tag_reg.re       = reg2hw.tag_601.re;
  assign rcache_line[2][89].status_reg.status = reg2hw.status_601.q;//status_reg_t'(reg2hw.status_601.q);
  assign rcache_line[2][89].status_reg.qe    = reg2hw.status_601.qe;
  assign rcache_line[2][89].status_reg.re    = reg2hw.status_601.re;


  assign rcache_line[2][90].tag_reg.tag      = reg2hw.tag_602.q;
  assign rcache_line[2][90].tag_reg.qe       = reg2hw.tag_602.qe;
  assign rcache_line[2][90].tag_reg.re       = reg2hw.tag_602.re;
  assign rcache_line[2][90].status_reg.status = reg2hw.status_602.q;//status_reg_t'(reg2hw.status_602.q);
  assign rcache_line[2][90].status_reg.qe    = reg2hw.status_602.qe;
  assign rcache_line[2][90].status_reg.re    = reg2hw.status_602.re;


  assign rcache_line[2][91].tag_reg.tag      = reg2hw.tag_603.q;
  assign rcache_line[2][91].tag_reg.qe       = reg2hw.tag_603.qe;
  assign rcache_line[2][91].tag_reg.re       = reg2hw.tag_603.re;
  assign rcache_line[2][91].status_reg.status = reg2hw.status_603.q;//status_reg_t'(reg2hw.status_603.q);
  assign rcache_line[2][91].status_reg.qe    = reg2hw.status_603.qe;
  assign rcache_line[2][91].status_reg.re    = reg2hw.status_603.re;


  assign rcache_line[2][92].tag_reg.tag      = reg2hw.tag_604.q;
  assign rcache_line[2][92].tag_reg.qe       = reg2hw.tag_604.qe;
  assign rcache_line[2][92].tag_reg.re       = reg2hw.tag_604.re;
  assign rcache_line[2][92].status_reg.status = reg2hw.status_604.q;//status_reg_t'(reg2hw.status_604.q);
  assign rcache_line[2][92].status_reg.qe    = reg2hw.status_604.qe;
  assign rcache_line[2][92].status_reg.re    = reg2hw.status_604.re;


  assign rcache_line[2][93].tag_reg.tag      = reg2hw.tag_605.q;
  assign rcache_line[2][93].tag_reg.qe       = reg2hw.tag_605.qe;
  assign rcache_line[2][93].tag_reg.re       = reg2hw.tag_605.re;
  assign rcache_line[2][93].status_reg.status = reg2hw.status_605.q;//status_reg_t'(reg2hw.status_605.q);
  assign rcache_line[2][93].status_reg.qe    = reg2hw.status_605.qe;
  assign rcache_line[2][93].status_reg.re    = reg2hw.status_605.re;


  assign rcache_line[2][94].tag_reg.tag      = reg2hw.tag_606.q;
  assign rcache_line[2][94].tag_reg.qe       = reg2hw.tag_606.qe;
  assign rcache_line[2][94].tag_reg.re       = reg2hw.tag_606.re;
  assign rcache_line[2][94].status_reg.status = reg2hw.status_606.q;//status_reg_t'(reg2hw.status_606.q);
  assign rcache_line[2][94].status_reg.qe    = reg2hw.status_606.qe;
  assign rcache_line[2][94].status_reg.re    = reg2hw.status_606.re;


  assign rcache_line[2][95].tag_reg.tag      = reg2hw.tag_607.q;
  assign rcache_line[2][95].tag_reg.qe       = reg2hw.tag_607.qe;
  assign rcache_line[2][95].tag_reg.re       = reg2hw.tag_607.re;
  assign rcache_line[2][95].status_reg.status = reg2hw.status_607.q;//status_reg_t'(reg2hw.status_607.q);
  assign rcache_line[2][95].status_reg.qe    = reg2hw.status_607.qe;
  assign rcache_line[2][95].status_reg.re    = reg2hw.status_607.re;


  assign rcache_line[2][96].tag_reg.tag      = reg2hw.tag_608.q;
  assign rcache_line[2][96].tag_reg.qe       = reg2hw.tag_608.qe;
  assign rcache_line[2][96].tag_reg.re       = reg2hw.tag_608.re;
  assign rcache_line[2][96].status_reg.status = reg2hw.status_608.q;//status_reg_t'(reg2hw.status_608.q);
  assign rcache_line[2][96].status_reg.qe    = reg2hw.status_608.qe;
  assign rcache_line[2][96].status_reg.re    = reg2hw.status_608.re;


  assign rcache_line[2][97].tag_reg.tag      = reg2hw.tag_609.q;
  assign rcache_line[2][97].tag_reg.qe       = reg2hw.tag_609.qe;
  assign rcache_line[2][97].tag_reg.re       = reg2hw.tag_609.re;
  assign rcache_line[2][97].status_reg.status = reg2hw.status_609.q;//status_reg_t'(reg2hw.status_609.q);
  assign rcache_line[2][97].status_reg.qe    = reg2hw.status_609.qe;
  assign rcache_line[2][97].status_reg.re    = reg2hw.status_609.re;


  assign rcache_line[2][98].tag_reg.tag      = reg2hw.tag_610.q;
  assign rcache_line[2][98].tag_reg.qe       = reg2hw.tag_610.qe;
  assign rcache_line[2][98].tag_reg.re       = reg2hw.tag_610.re;
  assign rcache_line[2][98].status_reg.status = reg2hw.status_610.q;//status_reg_t'(reg2hw.status_610.q);
  assign rcache_line[2][98].status_reg.qe    = reg2hw.status_610.qe;
  assign rcache_line[2][98].status_reg.re    = reg2hw.status_610.re;


  assign rcache_line[2][99].tag_reg.tag      = reg2hw.tag_611.q;
  assign rcache_line[2][99].tag_reg.qe       = reg2hw.tag_611.qe;
  assign rcache_line[2][99].tag_reg.re       = reg2hw.tag_611.re;
  assign rcache_line[2][99].status_reg.status = reg2hw.status_611.q;//status_reg_t'(reg2hw.status_611.q);
  assign rcache_line[2][99].status_reg.qe    = reg2hw.status_611.qe;
  assign rcache_line[2][99].status_reg.re    = reg2hw.status_611.re;


  assign rcache_line[2][100].tag_reg.tag      = reg2hw.tag_612.q;
  assign rcache_line[2][100].tag_reg.qe       = reg2hw.tag_612.qe;
  assign rcache_line[2][100].tag_reg.re       = reg2hw.tag_612.re;
  assign rcache_line[2][100].status_reg.status = reg2hw.status_612.q;//status_reg_t'(reg2hw.status_612.q);
  assign rcache_line[2][100].status_reg.qe    = reg2hw.status_612.qe;
  assign rcache_line[2][100].status_reg.re    = reg2hw.status_612.re;


  assign rcache_line[2][101].tag_reg.tag      = reg2hw.tag_613.q;
  assign rcache_line[2][101].tag_reg.qe       = reg2hw.tag_613.qe;
  assign rcache_line[2][101].tag_reg.re       = reg2hw.tag_613.re;
  assign rcache_line[2][101].status_reg.status = reg2hw.status_613.q;//status_reg_t'(reg2hw.status_613.q);
  assign rcache_line[2][101].status_reg.qe    = reg2hw.status_613.qe;
  assign rcache_line[2][101].status_reg.re    = reg2hw.status_613.re;


  assign rcache_line[2][102].tag_reg.tag      = reg2hw.tag_614.q;
  assign rcache_line[2][102].tag_reg.qe       = reg2hw.tag_614.qe;
  assign rcache_line[2][102].tag_reg.re       = reg2hw.tag_614.re;
  assign rcache_line[2][102].status_reg.status = reg2hw.status_614.q;//status_reg_t'(reg2hw.status_614.q);
  assign rcache_line[2][102].status_reg.qe    = reg2hw.status_614.qe;
  assign rcache_line[2][102].status_reg.re    = reg2hw.status_614.re;


  assign rcache_line[2][103].tag_reg.tag      = reg2hw.tag_615.q;
  assign rcache_line[2][103].tag_reg.qe       = reg2hw.tag_615.qe;
  assign rcache_line[2][103].tag_reg.re       = reg2hw.tag_615.re;
  assign rcache_line[2][103].status_reg.status = reg2hw.status_615.q;//status_reg_t'(reg2hw.status_615.q);
  assign rcache_line[2][103].status_reg.qe    = reg2hw.status_615.qe;
  assign rcache_line[2][103].status_reg.re    = reg2hw.status_615.re;


  assign rcache_line[2][104].tag_reg.tag      = reg2hw.tag_616.q;
  assign rcache_line[2][104].tag_reg.qe       = reg2hw.tag_616.qe;
  assign rcache_line[2][104].tag_reg.re       = reg2hw.tag_616.re;
  assign rcache_line[2][104].status_reg.status = reg2hw.status_616.q;//status_reg_t'(reg2hw.status_616.q);
  assign rcache_line[2][104].status_reg.qe    = reg2hw.status_616.qe;
  assign rcache_line[2][104].status_reg.re    = reg2hw.status_616.re;


  assign rcache_line[2][105].tag_reg.tag      = reg2hw.tag_617.q;
  assign rcache_line[2][105].tag_reg.qe       = reg2hw.tag_617.qe;
  assign rcache_line[2][105].tag_reg.re       = reg2hw.tag_617.re;
  assign rcache_line[2][105].status_reg.status = reg2hw.status_617.q;//status_reg_t'(reg2hw.status_617.q);
  assign rcache_line[2][105].status_reg.qe    = reg2hw.status_617.qe;
  assign rcache_line[2][105].status_reg.re    = reg2hw.status_617.re;


  assign rcache_line[2][106].tag_reg.tag      = reg2hw.tag_618.q;
  assign rcache_line[2][106].tag_reg.qe       = reg2hw.tag_618.qe;
  assign rcache_line[2][106].tag_reg.re       = reg2hw.tag_618.re;
  assign rcache_line[2][106].status_reg.status = reg2hw.status_618.q;//status_reg_t'(reg2hw.status_618.q);
  assign rcache_line[2][106].status_reg.qe    = reg2hw.status_618.qe;
  assign rcache_line[2][106].status_reg.re    = reg2hw.status_618.re;


  assign rcache_line[2][107].tag_reg.tag      = reg2hw.tag_619.q;
  assign rcache_line[2][107].tag_reg.qe       = reg2hw.tag_619.qe;
  assign rcache_line[2][107].tag_reg.re       = reg2hw.tag_619.re;
  assign rcache_line[2][107].status_reg.status = reg2hw.status_619.q;//status_reg_t'(reg2hw.status_619.q);
  assign rcache_line[2][107].status_reg.qe    = reg2hw.status_619.qe;
  assign rcache_line[2][107].status_reg.re    = reg2hw.status_619.re;


  assign rcache_line[2][108].tag_reg.tag      = reg2hw.tag_620.q;
  assign rcache_line[2][108].tag_reg.qe       = reg2hw.tag_620.qe;
  assign rcache_line[2][108].tag_reg.re       = reg2hw.tag_620.re;
  assign rcache_line[2][108].status_reg.status = reg2hw.status_620.q;//status_reg_t'(reg2hw.status_620.q);
  assign rcache_line[2][108].status_reg.qe    = reg2hw.status_620.qe;
  assign rcache_line[2][108].status_reg.re    = reg2hw.status_620.re;


  assign rcache_line[2][109].tag_reg.tag      = reg2hw.tag_621.q;
  assign rcache_line[2][109].tag_reg.qe       = reg2hw.tag_621.qe;
  assign rcache_line[2][109].tag_reg.re       = reg2hw.tag_621.re;
  assign rcache_line[2][109].status_reg.status = reg2hw.status_621.q;//status_reg_t'(reg2hw.status_621.q);
  assign rcache_line[2][109].status_reg.qe    = reg2hw.status_621.qe;
  assign rcache_line[2][109].status_reg.re    = reg2hw.status_621.re;


  assign rcache_line[2][110].tag_reg.tag      = reg2hw.tag_622.q;
  assign rcache_line[2][110].tag_reg.qe       = reg2hw.tag_622.qe;
  assign rcache_line[2][110].tag_reg.re       = reg2hw.tag_622.re;
  assign rcache_line[2][110].status_reg.status = reg2hw.status_622.q;//status_reg_t'(reg2hw.status_622.q);
  assign rcache_line[2][110].status_reg.qe    = reg2hw.status_622.qe;
  assign rcache_line[2][110].status_reg.re    = reg2hw.status_622.re;


  assign rcache_line[2][111].tag_reg.tag      = reg2hw.tag_623.q;
  assign rcache_line[2][111].tag_reg.qe       = reg2hw.tag_623.qe;
  assign rcache_line[2][111].tag_reg.re       = reg2hw.tag_623.re;
  assign rcache_line[2][111].status_reg.status = reg2hw.status_623.q;//status_reg_t'(reg2hw.status_623.q);
  assign rcache_line[2][111].status_reg.qe    = reg2hw.status_623.qe;
  assign rcache_line[2][111].status_reg.re    = reg2hw.status_623.re;


  assign rcache_line[2][112].tag_reg.tag      = reg2hw.tag_624.q;
  assign rcache_line[2][112].tag_reg.qe       = reg2hw.tag_624.qe;
  assign rcache_line[2][112].tag_reg.re       = reg2hw.tag_624.re;
  assign rcache_line[2][112].status_reg.status = reg2hw.status_624.q;//status_reg_t'(reg2hw.status_624.q);
  assign rcache_line[2][112].status_reg.qe    = reg2hw.status_624.qe;
  assign rcache_line[2][112].status_reg.re    = reg2hw.status_624.re;


  assign rcache_line[2][113].tag_reg.tag      = reg2hw.tag_625.q;
  assign rcache_line[2][113].tag_reg.qe       = reg2hw.tag_625.qe;
  assign rcache_line[2][113].tag_reg.re       = reg2hw.tag_625.re;
  assign rcache_line[2][113].status_reg.status = reg2hw.status_625.q;//status_reg_t'(reg2hw.status_625.q);
  assign rcache_line[2][113].status_reg.qe    = reg2hw.status_625.qe;
  assign rcache_line[2][113].status_reg.re    = reg2hw.status_625.re;


  assign rcache_line[2][114].tag_reg.tag      = reg2hw.tag_626.q;
  assign rcache_line[2][114].tag_reg.qe       = reg2hw.tag_626.qe;
  assign rcache_line[2][114].tag_reg.re       = reg2hw.tag_626.re;
  assign rcache_line[2][114].status_reg.status = reg2hw.status_626.q;//status_reg_t'(reg2hw.status_626.q);
  assign rcache_line[2][114].status_reg.qe    = reg2hw.status_626.qe;
  assign rcache_line[2][114].status_reg.re    = reg2hw.status_626.re;


  assign rcache_line[2][115].tag_reg.tag      = reg2hw.tag_627.q;
  assign rcache_line[2][115].tag_reg.qe       = reg2hw.tag_627.qe;
  assign rcache_line[2][115].tag_reg.re       = reg2hw.tag_627.re;
  assign rcache_line[2][115].status_reg.status = reg2hw.status_627.q;//status_reg_t'(reg2hw.status_627.q);
  assign rcache_line[2][115].status_reg.qe    = reg2hw.status_627.qe;
  assign rcache_line[2][115].status_reg.re    = reg2hw.status_627.re;


  assign rcache_line[2][116].tag_reg.tag      = reg2hw.tag_628.q;
  assign rcache_line[2][116].tag_reg.qe       = reg2hw.tag_628.qe;
  assign rcache_line[2][116].tag_reg.re       = reg2hw.tag_628.re;
  assign rcache_line[2][116].status_reg.status = reg2hw.status_628.q;//status_reg_t'(reg2hw.status_628.q);
  assign rcache_line[2][116].status_reg.qe    = reg2hw.status_628.qe;
  assign rcache_line[2][116].status_reg.re    = reg2hw.status_628.re;


  assign rcache_line[2][117].tag_reg.tag      = reg2hw.tag_629.q;
  assign rcache_line[2][117].tag_reg.qe       = reg2hw.tag_629.qe;
  assign rcache_line[2][117].tag_reg.re       = reg2hw.tag_629.re;
  assign rcache_line[2][117].status_reg.status = reg2hw.status_629.q;//status_reg_t'(reg2hw.status_629.q);
  assign rcache_line[2][117].status_reg.qe    = reg2hw.status_629.qe;
  assign rcache_line[2][117].status_reg.re    = reg2hw.status_629.re;


  assign rcache_line[2][118].tag_reg.tag      = reg2hw.tag_630.q;
  assign rcache_line[2][118].tag_reg.qe       = reg2hw.tag_630.qe;
  assign rcache_line[2][118].tag_reg.re       = reg2hw.tag_630.re;
  assign rcache_line[2][118].status_reg.status = reg2hw.status_630.q;//status_reg_t'(reg2hw.status_630.q);
  assign rcache_line[2][118].status_reg.qe    = reg2hw.status_630.qe;
  assign rcache_line[2][118].status_reg.re    = reg2hw.status_630.re;


  assign rcache_line[2][119].tag_reg.tag      = reg2hw.tag_631.q;
  assign rcache_line[2][119].tag_reg.qe       = reg2hw.tag_631.qe;
  assign rcache_line[2][119].tag_reg.re       = reg2hw.tag_631.re;
  assign rcache_line[2][119].status_reg.status = reg2hw.status_631.q;//status_reg_t'(reg2hw.status_631.q);
  assign rcache_line[2][119].status_reg.qe    = reg2hw.status_631.qe;
  assign rcache_line[2][119].status_reg.re    = reg2hw.status_631.re;


  assign rcache_line[2][120].tag_reg.tag      = reg2hw.tag_632.q;
  assign rcache_line[2][120].tag_reg.qe       = reg2hw.tag_632.qe;
  assign rcache_line[2][120].tag_reg.re       = reg2hw.tag_632.re;
  assign rcache_line[2][120].status_reg.status = reg2hw.status_632.q;//status_reg_t'(reg2hw.status_632.q);
  assign rcache_line[2][120].status_reg.qe    = reg2hw.status_632.qe;
  assign rcache_line[2][120].status_reg.re    = reg2hw.status_632.re;


  assign rcache_line[2][121].tag_reg.tag      = reg2hw.tag_633.q;
  assign rcache_line[2][121].tag_reg.qe       = reg2hw.tag_633.qe;
  assign rcache_line[2][121].tag_reg.re       = reg2hw.tag_633.re;
  assign rcache_line[2][121].status_reg.status = reg2hw.status_633.q;//status_reg_t'(reg2hw.status_633.q);
  assign rcache_line[2][121].status_reg.qe    = reg2hw.status_633.qe;
  assign rcache_line[2][121].status_reg.re    = reg2hw.status_633.re;


  assign rcache_line[2][122].tag_reg.tag      = reg2hw.tag_634.q;
  assign rcache_line[2][122].tag_reg.qe       = reg2hw.tag_634.qe;
  assign rcache_line[2][122].tag_reg.re       = reg2hw.tag_634.re;
  assign rcache_line[2][122].status_reg.status = reg2hw.status_634.q;//status_reg_t'(reg2hw.status_634.q);
  assign rcache_line[2][122].status_reg.qe    = reg2hw.status_634.qe;
  assign rcache_line[2][122].status_reg.re    = reg2hw.status_634.re;


  assign rcache_line[2][123].tag_reg.tag      = reg2hw.tag_635.q;
  assign rcache_line[2][123].tag_reg.qe       = reg2hw.tag_635.qe;
  assign rcache_line[2][123].tag_reg.re       = reg2hw.tag_635.re;
  assign rcache_line[2][123].status_reg.status = reg2hw.status_635.q;//status_reg_t'(reg2hw.status_635.q);
  assign rcache_line[2][123].status_reg.qe    = reg2hw.status_635.qe;
  assign rcache_line[2][123].status_reg.re    = reg2hw.status_635.re;


  assign rcache_line[2][124].tag_reg.tag      = reg2hw.tag_636.q;
  assign rcache_line[2][124].tag_reg.qe       = reg2hw.tag_636.qe;
  assign rcache_line[2][124].tag_reg.re       = reg2hw.tag_636.re;
  assign rcache_line[2][124].status_reg.status = reg2hw.status_636.q;//status_reg_t'(reg2hw.status_636.q);
  assign rcache_line[2][124].status_reg.qe    = reg2hw.status_636.qe;
  assign rcache_line[2][124].status_reg.re    = reg2hw.status_636.re;


  assign rcache_line[2][125].tag_reg.tag      = reg2hw.tag_637.q;
  assign rcache_line[2][125].tag_reg.qe       = reg2hw.tag_637.qe;
  assign rcache_line[2][125].tag_reg.re       = reg2hw.tag_637.re;
  assign rcache_line[2][125].status_reg.status = reg2hw.status_637.q;//status_reg_t'(reg2hw.status_637.q);
  assign rcache_line[2][125].status_reg.qe    = reg2hw.status_637.qe;
  assign rcache_line[2][125].status_reg.re    = reg2hw.status_637.re;


  assign rcache_line[2][126].tag_reg.tag      = reg2hw.tag_638.q;
  assign rcache_line[2][126].tag_reg.qe       = reg2hw.tag_638.qe;
  assign rcache_line[2][126].tag_reg.re       = reg2hw.tag_638.re;
  assign rcache_line[2][126].status_reg.status = reg2hw.status_638.q;//status_reg_t'(reg2hw.status_638.q);
  assign rcache_line[2][126].status_reg.qe    = reg2hw.status_638.qe;
  assign rcache_line[2][126].status_reg.re    = reg2hw.status_638.re;


  assign rcache_line[2][127].tag_reg.tag      = reg2hw.tag_639.q;
  assign rcache_line[2][127].tag_reg.qe       = reg2hw.tag_639.qe;
  assign rcache_line[2][127].tag_reg.re       = reg2hw.tag_639.re;
  assign rcache_line[2][127].status_reg.status = reg2hw.status_639.q;//status_reg_t'(reg2hw.status_639.q);
  assign rcache_line[2][127].status_reg.qe    = reg2hw.status_639.qe;
  assign rcache_line[2][127].status_reg.re    = reg2hw.status_639.re;


  assign rcache_line[2][128].tag_reg.tag      = reg2hw.tag_640.q;
  assign rcache_line[2][128].tag_reg.qe       = reg2hw.tag_640.qe;
  assign rcache_line[2][128].tag_reg.re       = reg2hw.tag_640.re;
  assign rcache_line[2][128].status_reg.status = reg2hw.status_640.q;//status_reg_t'(reg2hw.status_640.q);
  assign rcache_line[2][128].status_reg.qe    = reg2hw.status_640.qe;
  assign rcache_line[2][128].status_reg.re    = reg2hw.status_640.re;


  assign rcache_line[2][129].tag_reg.tag      = reg2hw.tag_641.q;
  assign rcache_line[2][129].tag_reg.qe       = reg2hw.tag_641.qe;
  assign rcache_line[2][129].tag_reg.re       = reg2hw.tag_641.re;
  assign rcache_line[2][129].status_reg.status = reg2hw.status_641.q;//status_reg_t'(reg2hw.status_641.q);
  assign rcache_line[2][129].status_reg.qe    = reg2hw.status_641.qe;
  assign rcache_line[2][129].status_reg.re    = reg2hw.status_641.re;


  assign rcache_line[2][130].tag_reg.tag      = reg2hw.tag_642.q;
  assign rcache_line[2][130].tag_reg.qe       = reg2hw.tag_642.qe;
  assign rcache_line[2][130].tag_reg.re       = reg2hw.tag_642.re;
  assign rcache_line[2][130].status_reg.status = reg2hw.status_642.q;//status_reg_t'(reg2hw.status_642.q);
  assign rcache_line[2][130].status_reg.qe    = reg2hw.status_642.qe;
  assign rcache_line[2][130].status_reg.re    = reg2hw.status_642.re;


  assign rcache_line[2][131].tag_reg.tag      = reg2hw.tag_643.q;
  assign rcache_line[2][131].tag_reg.qe       = reg2hw.tag_643.qe;
  assign rcache_line[2][131].tag_reg.re       = reg2hw.tag_643.re;
  assign rcache_line[2][131].status_reg.status = reg2hw.status_643.q;//status_reg_t'(reg2hw.status_643.q);
  assign rcache_line[2][131].status_reg.qe    = reg2hw.status_643.qe;
  assign rcache_line[2][131].status_reg.re    = reg2hw.status_643.re;


  assign rcache_line[2][132].tag_reg.tag      = reg2hw.tag_644.q;
  assign rcache_line[2][132].tag_reg.qe       = reg2hw.tag_644.qe;
  assign rcache_line[2][132].tag_reg.re       = reg2hw.tag_644.re;
  assign rcache_line[2][132].status_reg.status = reg2hw.status_644.q;//status_reg_t'(reg2hw.status_644.q);
  assign rcache_line[2][132].status_reg.qe    = reg2hw.status_644.qe;
  assign rcache_line[2][132].status_reg.re    = reg2hw.status_644.re;


  assign rcache_line[2][133].tag_reg.tag      = reg2hw.tag_645.q;
  assign rcache_line[2][133].tag_reg.qe       = reg2hw.tag_645.qe;
  assign rcache_line[2][133].tag_reg.re       = reg2hw.tag_645.re;
  assign rcache_line[2][133].status_reg.status = reg2hw.status_645.q;//status_reg_t'(reg2hw.status_645.q);
  assign rcache_line[2][133].status_reg.qe    = reg2hw.status_645.qe;
  assign rcache_line[2][133].status_reg.re    = reg2hw.status_645.re;


  assign rcache_line[2][134].tag_reg.tag      = reg2hw.tag_646.q;
  assign rcache_line[2][134].tag_reg.qe       = reg2hw.tag_646.qe;
  assign rcache_line[2][134].tag_reg.re       = reg2hw.tag_646.re;
  assign rcache_line[2][134].status_reg.status = reg2hw.status_646.q;//status_reg_t'(reg2hw.status_646.q);
  assign rcache_line[2][134].status_reg.qe    = reg2hw.status_646.qe;
  assign rcache_line[2][134].status_reg.re    = reg2hw.status_646.re;


  assign rcache_line[2][135].tag_reg.tag      = reg2hw.tag_647.q;
  assign rcache_line[2][135].tag_reg.qe       = reg2hw.tag_647.qe;
  assign rcache_line[2][135].tag_reg.re       = reg2hw.tag_647.re;
  assign rcache_line[2][135].status_reg.status = reg2hw.status_647.q;//status_reg_t'(reg2hw.status_647.q);
  assign rcache_line[2][135].status_reg.qe    = reg2hw.status_647.qe;
  assign rcache_line[2][135].status_reg.re    = reg2hw.status_647.re;


  assign rcache_line[2][136].tag_reg.tag      = reg2hw.tag_648.q;
  assign rcache_line[2][136].tag_reg.qe       = reg2hw.tag_648.qe;
  assign rcache_line[2][136].tag_reg.re       = reg2hw.tag_648.re;
  assign rcache_line[2][136].status_reg.status = reg2hw.status_648.q;//status_reg_t'(reg2hw.status_648.q);
  assign rcache_line[2][136].status_reg.qe    = reg2hw.status_648.qe;
  assign rcache_line[2][136].status_reg.re    = reg2hw.status_648.re;


  assign rcache_line[2][137].tag_reg.tag      = reg2hw.tag_649.q;
  assign rcache_line[2][137].tag_reg.qe       = reg2hw.tag_649.qe;
  assign rcache_line[2][137].tag_reg.re       = reg2hw.tag_649.re;
  assign rcache_line[2][137].status_reg.status = reg2hw.status_649.q;//status_reg_t'(reg2hw.status_649.q);
  assign rcache_line[2][137].status_reg.qe    = reg2hw.status_649.qe;
  assign rcache_line[2][137].status_reg.re    = reg2hw.status_649.re;


  assign rcache_line[2][138].tag_reg.tag      = reg2hw.tag_650.q;
  assign rcache_line[2][138].tag_reg.qe       = reg2hw.tag_650.qe;
  assign rcache_line[2][138].tag_reg.re       = reg2hw.tag_650.re;
  assign rcache_line[2][138].status_reg.status = reg2hw.status_650.q;//status_reg_t'(reg2hw.status_650.q);
  assign rcache_line[2][138].status_reg.qe    = reg2hw.status_650.qe;
  assign rcache_line[2][138].status_reg.re    = reg2hw.status_650.re;


  assign rcache_line[2][139].tag_reg.tag      = reg2hw.tag_651.q;
  assign rcache_line[2][139].tag_reg.qe       = reg2hw.tag_651.qe;
  assign rcache_line[2][139].tag_reg.re       = reg2hw.tag_651.re;
  assign rcache_line[2][139].status_reg.status = reg2hw.status_651.q;//status_reg_t'(reg2hw.status_651.q);
  assign rcache_line[2][139].status_reg.qe    = reg2hw.status_651.qe;
  assign rcache_line[2][139].status_reg.re    = reg2hw.status_651.re;


  assign rcache_line[2][140].tag_reg.tag      = reg2hw.tag_652.q;
  assign rcache_line[2][140].tag_reg.qe       = reg2hw.tag_652.qe;
  assign rcache_line[2][140].tag_reg.re       = reg2hw.tag_652.re;
  assign rcache_line[2][140].status_reg.status = reg2hw.status_652.q;//status_reg_t'(reg2hw.status_652.q);
  assign rcache_line[2][140].status_reg.qe    = reg2hw.status_652.qe;
  assign rcache_line[2][140].status_reg.re    = reg2hw.status_652.re;


  assign rcache_line[2][141].tag_reg.tag      = reg2hw.tag_653.q;
  assign rcache_line[2][141].tag_reg.qe       = reg2hw.tag_653.qe;
  assign rcache_line[2][141].tag_reg.re       = reg2hw.tag_653.re;
  assign rcache_line[2][141].status_reg.status = reg2hw.status_653.q;//status_reg_t'(reg2hw.status_653.q);
  assign rcache_line[2][141].status_reg.qe    = reg2hw.status_653.qe;
  assign rcache_line[2][141].status_reg.re    = reg2hw.status_653.re;


  assign rcache_line[2][142].tag_reg.tag      = reg2hw.tag_654.q;
  assign rcache_line[2][142].tag_reg.qe       = reg2hw.tag_654.qe;
  assign rcache_line[2][142].tag_reg.re       = reg2hw.tag_654.re;
  assign rcache_line[2][142].status_reg.status = reg2hw.status_654.q;//status_reg_t'(reg2hw.status_654.q);
  assign rcache_line[2][142].status_reg.qe    = reg2hw.status_654.qe;
  assign rcache_line[2][142].status_reg.re    = reg2hw.status_654.re;


  assign rcache_line[2][143].tag_reg.tag      = reg2hw.tag_655.q;
  assign rcache_line[2][143].tag_reg.qe       = reg2hw.tag_655.qe;
  assign rcache_line[2][143].tag_reg.re       = reg2hw.tag_655.re;
  assign rcache_line[2][143].status_reg.status = reg2hw.status_655.q;//status_reg_t'(reg2hw.status_655.q);
  assign rcache_line[2][143].status_reg.qe    = reg2hw.status_655.qe;
  assign rcache_line[2][143].status_reg.re    = reg2hw.status_655.re;


  assign rcache_line[2][144].tag_reg.tag      = reg2hw.tag_656.q;
  assign rcache_line[2][144].tag_reg.qe       = reg2hw.tag_656.qe;
  assign rcache_line[2][144].tag_reg.re       = reg2hw.tag_656.re;
  assign rcache_line[2][144].status_reg.status = reg2hw.status_656.q;//status_reg_t'(reg2hw.status_656.q);
  assign rcache_line[2][144].status_reg.qe    = reg2hw.status_656.qe;
  assign rcache_line[2][144].status_reg.re    = reg2hw.status_656.re;


  assign rcache_line[2][145].tag_reg.tag      = reg2hw.tag_657.q;
  assign rcache_line[2][145].tag_reg.qe       = reg2hw.tag_657.qe;
  assign rcache_line[2][145].tag_reg.re       = reg2hw.tag_657.re;
  assign rcache_line[2][145].status_reg.status = reg2hw.status_657.q;//status_reg_t'(reg2hw.status_657.q);
  assign rcache_line[2][145].status_reg.qe    = reg2hw.status_657.qe;
  assign rcache_line[2][145].status_reg.re    = reg2hw.status_657.re;


  assign rcache_line[2][146].tag_reg.tag      = reg2hw.tag_658.q;
  assign rcache_line[2][146].tag_reg.qe       = reg2hw.tag_658.qe;
  assign rcache_line[2][146].tag_reg.re       = reg2hw.tag_658.re;
  assign rcache_line[2][146].status_reg.status = reg2hw.status_658.q;//status_reg_t'(reg2hw.status_658.q);
  assign rcache_line[2][146].status_reg.qe    = reg2hw.status_658.qe;
  assign rcache_line[2][146].status_reg.re    = reg2hw.status_658.re;


  assign rcache_line[2][147].tag_reg.tag      = reg2hw.tag_659.q;
  assign rcache_line[2][147].tag_reg.qe       = reg2hw.tag_659.qe;
  assign rcache_line[2][147].tag_reg.re       = reg2hw.tag_659.re;
  assign rcache_line[2][147].status_reg.status = reg2hw.status_659.q;//status_reg_t'(reg2hw.status_659.q);
  assign rcache_line[2][147].status_reg.qe    = reg2hw.status_659.qe;
  assign rcache_line[2][147].status_reg.re    = reg2hw.status_659.re;


  assign rcache_line[2][148].tag_reg.tag      = reg2hw.tag_660.q;
  assign rcache_line[2][148].tag_reg.qe       = reg2hw.tag_660.qe;
  assign rcache_line[2][148].tag_reg.re       = reg2hw.tag_660.re;
  assign rcache_line[2][148].status_reg.status = reg2hw.status_660.q;//status_reg_t'(reg2hw.status_660.q);
  assign rcache_line[2][148].status_reg.qe    = reg2hw.status_660.qe;
  assign rcache_line[2][148].status_reg.re    = reg2hw.status_660.re;


  assign rcache_line[2][149].tag_reg.tag      = reg2hw.tag_661.q;
  assign rcache_line[2][149].tag_reg.qe       = reg2hw.tag_661.qe;
  assign rcache_line[2][149].tag_reg.re       = reg2hw.tag_661.re;
  assign rcache_line[2][149].status_reg.status = reg2hw.status_661.q;//status_reg_t'(reg2hw.status_661.q);
  assign rcache_line[2][149].status_reg.qe    = reg2hw.status_661.qe;
  assign rcache_line[2][149].status_reg.re    = reg2hw.status_661.re;


  assign rcache_line[2][150].tag_reg.tag      = reg2hw.tag_662.q;
  assign rcache_line[2][150].tag_reg.qe       = reg2hw.tag_662.qe;
  assign rcache_line[2][150].tag_reg.re       = reg2hw.tag_662.re;
  assign rcache_line[2][150].status_reg.status = reg2hw.status_662.q;//status_reg_t'(reg2hw.status_662.q);
  assign rcache_line[2][150].status_reg.qe    = reg2hw.status_662.qe;
  assign rcache_line[2][150].status_reg.re    = reg2hw.status_662.re;


  assign rcache_line[2][151].tag_reg.tag      = reg2hw.tag_663.q;
  assign rcache_line[2][151].tag_reg.qe       = reg2hw.tag_663.qe;
  assign rcache_line[2][151].tag_reg.re       = reg2hw.tag_663.re;
  assign rcache_line[2][151].status_reg.status = reg2hw.status_663.q;//status_reg_t'(reg2hw.status_663.q);
  assign rcache_line[2][151].status_reg.qe    = reg2hw.status_663.qe;
  assign rcache_line[2][151].status_reg.re    = reg2hw.status_663.re;


  assign rcache_line[2][152].tag_reg.tag      = reg2hw.tag_664.q;
  assign rcache_line[2][152].tag_reg.qe       = reg2hw.tag_664.qe;
  assign rcache_line[2][152].tag_reg.re       = reg2hw.tag_664.re;
  assign rcache_line[2][152].status_reg.status = reg2hw.status_664.q;//status_reg_t'(reg2hw.status_664.q);
  assign rcache_line[2][152].status_reg.qe    = reg2hw.status_664.qe;
  assign rcache_line[2][152].status_reg.re    = reg2hw.status_664.re;


  assign rcache_line[2][153].tag_reg.tag      = reg2hw.tag_665.q;
  assign rcache_line[2][153].tag_reg.qe       = reg2hw.tag_665.qe;
  assign rcache_line[2][153].tag_reg.re       = reg2hw.tag_665.re;
  assign rcache_line[2][153].status_reg.status = reg2hw.status_665.q;//status_reg_t'(reg2hw.status_665.q);
  assign rcache_line[2][153].status_reg.qe    = reg2hw.status_665.qe;
  assign rcache_line[2][153].status_reg.re    = reg2hw.status_665.re;


  assign rcache_line[2][154].tag_reg.tag      = reg2hw.tag_666.q;
  assign rcache_line[2][154].tag_reg.qe       = reg2hw.tag_666.qe;
  assign rcache_line[2][154].tag_reg.re       = reg2hw.tag_666.re;
  assign rcache_line[2][154].status_reg.status = reg2hw.status_666.q;//status_reg_t'(reg2hw.status_666.q);
  assign rcache_line[2][154].status_reg.qe    = reg2hw.status_666.qe;
  assign rcache_line[2][154].status_reg.re    = reg2hw.status_666.re;


  assign rcache_line[2][155].tag_reg.tag      = reg2hw.tag_667.q;
  assign rcache_line[2][155].tag_reg.qe       = reg2hw.tag_667.qe;
  assign rcache_line[2][155].tag_reg.re       = reg2hw.tag_667.re;
  assign rcache_line[2][155].status_reg.status = reg2hw.status_667.q;//status_reg_t'(reg2hw.status_667.q);
  assign rcache_line[2][155].status_reg.qe    = reg2hw.status_667.qe;
  assign rcache_line[2][155].status_reg.re    = reg2hw.status_667.re;


  assign rcache_line[2][156].tag_reg.tag      = reg2hw.tag_668.q;
  assign rcache_line[2][156].tag_reg.qe       = reg2hw.tag_668.qe;
  assign rcache_line[2][156].tag_reg.re       = reg2hw.tag_668.re;
  assign rcache_line[2][156].status_reg.status = reg2hw.status_668.q;//status_reg_t'(reg2hw.status_668.q);
  assign rcache_line[2][156].status_reg.qe    = reg2hw.status_668.qe;
  assign rcache_line[2][156].status_reg.re    = reg2hw.status_668.re;


  assign rcache_line[2][157].tag_reg.tag      = reg2hw.tag_669.q;
  assign rcache_line[2][157].tag_reg.qe       = reg2hw.tag_669.qe;
  assign rcache_line[2][157].tag_reg.re       = reg2hw.tag_669.re;
  assign rcache_line[2][157].status_reg.status = reg2hw.status_669.q;//status_reg_t'(reg2hw.status_669.q);
  assign rcache_line[2][157].status_reg.qe    = reg2hw.status_669.qe;
  assign rcache_line[2][157].status_reg.re    = reg2hw.status_669.re;


  assign rcache_line[2][158].tag_reg.tag      = reg2hw.tag_670.q;
  assign rcache_line[2][158].tag_reg.qe       = reg2hw.tag_670.qe;
  assign rcache_line[2][158].tag_reg.re       = reg2hw.tag_670.re;
  assign rcache_line[2][158].status_reg.status = reg2hw.status_670.q;//status_reg_t'(reg2hw.status_670.q);
  assign rcache_line[2][158].status_reg.qe    = reg2hw.status_670.qe;
  assign rcache_line[2][158].status_reg.re    = reg2hw.status_670.re;


  assign rcache_line[2][159].tag_reg.tag      = reg2hw.tag_671.q;
  assign rcache_line[2][159].tag_reg.qe       = reg2hw.tag_671.qe;
  assign rcache_line[2][159].tag_reg.re       = reg2hw.tag_671.re;
  assign rcache_line[2][159].status_reg.status = reg2hw.status_671.q;//status_reg_t'(reg2hw.status_671.q);
  assign rcache_line[2][159].status_reg.qe    = reg2hw.status_671.qe;
  assign rcache_line[2][159].status_reg.re    = reg2hw.status_671.re;


  assign rcache_line[2][160].tag_reg.tag      = reg2hw.tag_672.q;
  assign rcache_line[2][160].tag_reg.qe       = reg2hw.tag_672.qe;
  assign rcache_line[2][160].tag_reg.re       = reg2hw.tag_672.re;
  assign rcache_line[2][160].status_reg.status = reg2hw.status_672.q;//status_reg_t'(reg2hw.status_672.q);
  assign rcache_line[2][160].status_reg.qe    = reg2hw.status_672.qe;
  assign rcache_line[2][160].status_reg.re    = reg2hw.status_672.re;


  assign rcache_line[2][161].tag_reg.tag      = reg2hw.tag_673.q;
  assign rcache_line[2][161].tag_reg.qe       = reg2hw.tag_673.qe;
  assign rcache_line[2][161].tag_reg.re       = reg2hw.tag_673.re;
  assign rcache_line[2][161].status_reg.status = reg2hw.status_673.q;//status_reg_t'(reg2hw.status_673.q);
  assign rcache_line[2][161].status_reg.qe    = reg2hw.status_673.qe;
  assign rcache_line[2][161].status_reg.re    = reg2hw.status_673.re;


  assign rcache_line[2][162].tag_reg.tag      = reg2hw.tag_674.q;
  assign rcache_line[2][162].tag_reg.qe       = reg2hw.tag_674.qe;
  assign rcache_line[2][162].tag_reg.re       = reg2hw.tag_674.re;
  assign rcache_line[2][162].status_reg.status = reg2hw.status_674.q;//status_reg_t'(reg2hw.status_674.q);
  assign rcache_line[2][162].status_reg.qe    = reg2hw.status_674.qe;
  assign rcache_line[2][162].status_reg.re    = reg2hw.status_674.re;


  assign rcache_line[2][163].tag_reg.tag      = reg2hw.tag_675.q;
  assign rcache_line[2][163].tag_reg.qe       = reg2hw.tag_675.qe;
  assign rcache_line[2][163].tag_reg.re       = reg2hw.tag_675.re;
  assign rcache_line[2][163].status_reg.status = reg2hw.status_675.q;//status_reg_t'(reg2hw.status_675.q);
  assign rcache_line[2][163].status_reg.qe    = reg2hw.status_675.qe;
  assign rcache_line[2][163].status_reg.re    = reg2hw.status_675.re;


  assign rcache_line[2][164].tag_reg.tag      = reg2hw.tag_676.q;
  assign rcache_line[2][164].tag_reg.qe       = reg2hw.tag_676.qe;
  assign rcache_line[2][164].tag_reg.re       = reg2hw.tag_676.re;
  assign rcache_line[2][164].status_reg.status = reg2hw.status_676.q;//status_reg_t'(reg2hw.status_676.q);
  assign rcache_line[2][164].status_reg.qe    = reg2hw.status_676.qe;
  assign rcache_line[2][164].status_reg.re    = reg2hw.status_676.re;


  assign rcache_line[2][165].tag_reg.tag      = reg2hw.tag_677.q;
  assign rcache_line[2][165].tag_reg.qe       = reg2hw.tag_677.qe;
  assign rcache_line[2][165].tag_reg.re       = reg2hw.tag_677.re;
  assign rcache_line[2][165].status_reg.status = reg2hw.status_677.q;//status_reg_t'(reg2hw.status_677.q);
  assign rcache_line[2][165].status_reg.qe    = reg2hw.status_677.qe;
  assign rcache_line[2][165].status_reg.re    = reg2hw.status_677.re;


  assign rcache_line[2][166].tag_reg.tag      = reg2hw.tag_678.q;
  assign rcache_line[2][166].tag_reg.qe       = reg2hw.tag_678.qe;
  assign rcache_line[2][166].tag_reg.re       = reg2hw.tag_678.re;
  assign rcache_line[2][166].status_reg.status = reg2hw.status_678.q;//status_reg_t'(reg2hw.status_678.q);
  assign rcache_line[2][166].status_reg.qe    = reg2hw.status_678.qe;
  assign rcache_line[2][166].status_reg.re    = reg2hw.status_678.re;


  assign rcache_line[2][167].tag_reg.tag      = reg2hw.tag_679.q;
  assign rcache_line[2][167].tag_reg.qe       = reg2hw.tag_679.qe;
  assign rcache_line[2][167].tag_reg.re       = reg2hw.tag_679.re;
  assign rcache_line[2][167].status_reg.status = reg2hw.status_679.q;//status_reg_t'(reg2hw.status_679.q);
  assign rcache_line[2][167].status_reg.qe    = reg2hw.status_679.qe;
  assign rcache_line[2][167].status_reg.re    = reg2hw.status_679.re;


  assign rcache_line[2][168].tag_reg.tag      = reg2hw.tag_680.q;
  assign rcache_line[2][168].tag_reg.qe       = reg2hw.tag_680.qe;
  assign rcache_line[2][168].tag_reg.re       = reg2hw.tag_680.re;
  assign rcache_line[2][168].status_reg.status = reg2hw.status_680.q;//status_reg_t'(reg2hw.status_680.q);
  assign rcache_line[2][168].status_reg.qe    = reg2hw.status_680.qe;
  assign rcache_line[2][168].status_reg.re    = reg2hw.status_680.re;


  assign rcache_line[2][169].tag_reg.tag      = reg2hw.tag_681.q;
  assign rcache_line[2][169].tag_reg.qe       = reg2hw.tag_681.qe;
  assign rcache_line[2][169].tag_reg.re       = reg2hw.tag_681.re;
  assign rcache_line[2][169].status_reg.status = reg2hw.status_681.q;//status_reg_t'(reg2hw.status_681.q);
  assign rcache_line[2][169].status_reg.qe    = reg2hw.status_681.qe;
  assign rcache_line[2][169].status_reg.re    = reg2hw.status_681.re;


  assign rcache_line[2][170].tag_reg.tag      = reg2hw.tag_682.q;
  assign rcache_line[2][170].tag_reg.qe       = reg2hw.tag_682.qe;
  assign rcache_line[2][170].tag_reg.re       = reg2hw.tag_682.re;
  assign rcache_line[2][170].status_reg.status = reg2hw.status_682.q;//status_reg_t'(reg2hw.status_682.q);
  assign rcache_line[2][170].status_reg.qe    = reg2hw.status_682.qe;
  assign rcache_line[2][170].status_reg.re    = reg2hw.status_682.re;


  assign rcache_line[2][171].tag_reg.tag      = reg2hw.tag_683.q;
  assign rcache_line[2][171].tag_reg.qe       = reg2hw.tag_683.qe;
  assign rcache_line[2][171].tag_reg.re       = reg2hw.tag_683.re;
  assign rcache_line[2][171].status_reg.status = reg2hw.status_683.q;//status_reg_t'(reg2hw.status_683.q);
  assign rcache_line[2][171].status_reg.qe    = reg2hw.status_683.qe;
  assign rcache_line[2][171].status_reg.re    = reg2hw.status_683.re;


  assign rcache_line[2][172].tag_reg.tag      = reg2hw.tag_684.q;
  assign rcache_line[2][172].tag_reg.qe       = reg2hw.tag_684.qe;
  assign rcache_line[2][172].tag_reg.re       = reg2hw.tag_684.re;
  assign rcache_line[2][172].status_reg.status = reg2hw.status_684.q;//status_reg_t'(reg2hw.status_684.q);
  assign rcache_line[2][172].status_reg.qe    = reg2hw.status_684.qe;
  assign rcache_line[2][172].status_reg.re    = reg2hw.status_684.re;


  assign rcache_line[2][173].tag_reg.tag      = reg2hw.tag_685.q;
  assign rcache_line[2][173].tag_reg.qe       = reg2hw.tag_685.qe;
  assign rcache_line[2][173].tag_reg.re       = reg2hw.tag_685.re;
  assign rcache_line[2][173].status_reg.status = reg2hw.status_685.q;//status_reg_t'(reg2hw.status_685.q);
  assign rcache_line[2][173].status_reg.qe    = reg2hw.status_685.qe;
  assign rcache_line[2][173].status_reg.re    = reg2hw.status_685.re;


  assign rcache_line[2][174].tag_reg.tag      = reg2hw.tag_686.q;
  assign rcache_line[2][174].tag_reg.qe       = reg2hw.tag_686.qe;
  assign rcache_line[2][174].tag_reg.re       = reg2hw.tag_686.re;
  assign rcache_line[2][174].status_reg.status = reg2hw.status_686.q;//status_reg_t'(reg2hw.status_686.q);
  assign rcache_line[2][174].status_reg.qe    = reg2hw.status_686.qe;
  assign rcache_line[2][174].status_reg.re    = reg2hw.status_686.re;


  assign rcache_line[2][175].tag_reg.tag      = reg2hw.tag_687.q;
  assign rcache_line[2][175].tag_reg.qe       = reg2hw.tag_687.qe;
  assign rcache_line[2][175].tag_reg.re       = reg2hw.tag_687.re;
  assign rcache_line[2][175].status_reg.status = reg2hw.status_687.q;//status_reg_t'(reg2hw.status_687.q);
  assign rcache_line[2][175].status_reg.qe    = reg2hw.status_687.qe;
  assign rcache_line[2][175].status_reg.re    = reg2hw.status_687.re;


  assign rcache_line[2][176].tag_reg.tag      = reg2hw.tag_688.q;
  assign rcache_line[2][176].tag_reg.qe       = reg2hw.tag_688.qe;
  assign rcache_line[2][176].tag_reg.re       = reg2hw.tag_688.re;
  assign rcache_line[2][176].status_reg.status = reg2hw.status_688.q;//status_reg_t'(reg2hw.status_688.q);
  assign rcache_line[2][176].status_reg.qe    = reg2hw.status_688.qe;
  assign rcache_line[2][176].status_reg.re    = reg2hw.status_688.re;


  assign rcache_line[2][177].tag_reg.tag      = reg2hw.tag_689.q;
  assign rcache_line[2][177].tag_reg.qe       = reg2hw.tag_689.qe;
  assign rcache_line[2][177].tag_reg.re       = reg2hw.tag_689.re;
  assign rcache_line[2][177].status_reg.status = reg2hw.status_689.q;//status_reg_t'(reg2hw.status_689.q);
  assign rcache_line[2][177].status_reg.qe    = reg2hw.status_689.qe;
  assign rcache_line[2][177].status_reg.re    = reg2hw.status_689.re;


  assign rcache_line[2][178].tag_reg.tag      = reg2hw.tag_690.q;
  assign rcache_line[2][178].tag_reg.qe       = reg2hw.tag_690.qe;
  assign rcache_line[2][178].tag_reg.re       = reg2hw.tag_690.re;
  assign rcache_line[2][178].status_reg.status = reg2hw.status_690.q;//status_reg_t'(reg2hw.status_690.q);
  assign rcache_line[2][178].status_reg.qe    = reg2hw.status_690.qe;
  assign rcache_line[2][178].status_reg.re    = reg2hw.status_690.re;


  assign rcache_line[2][179].tag_reg.tag      = reg2hw.tag_691.q;
  assign rcache_line[2][179].tag_reg.qe       = reg2hw.tag_691.qe;
  assign rcache_line[2][179].tag_reg.re       = reg2hw.tag_691.re;
  assign rcache_line[2][179].status_reg.status = reg2hw.status_691.q;//status_reg_t'(reg2hw.status_691.q);
  assign rcache_line[2][179].status_reg.qe    = reg2hw.status_691.qe;
  assign rcache_line[2][179].status_reg.re    = reg2hw.status_691.re;


  assign rcache_line[2][180].tag_reg.tag      = reg2hw.tag_692.q;
  assign rcache_line[2][180].tag_reg.qe       = reg2hw.tag_692.qe;
  assign rcache_line[2][180].tag_reg.re       = reg2hw.tag_692.re;
  assign rcache_line[2][180].status_reg.status = reg2hw.status_692.q;//status_reg_t'(reg2hw.status_692.q);
  assign rcache_line[2][180].status_reg.qe    = reg2hw.status_692.qe;
  assign rcache_line[2][180].status_reg.re    = reg2hw.status_692.re;


  assign rcache_line[2][181].tag_reg.tag      = reg2hw.tag_693.q;
  assign rcache_line[2][181].tag_reg.qe       = reg2hw.tag_693.qe;
  assign rcache_line[2][181].tag_reg.re       = reg2hw.tag_693.re;
  assign rcache_line[2][181].status_reg.status = reg2hw.status_693.q;//status_reg_t'(reg2hw.status_693.q);
  assign rcache_line[2][181].status_reg.qe    = reg2hw.status_693.qe;
  assign rcache_line[2][181].status_reg.re    = reg2hw.status_693.re;


  assign rcache_line[2][182].tag_reg.tag      = reg2hw.tag_694.q;
  assign rcache_line[2][182].tag_reg.qe       = reg2hw.tag_694.qe;
  assign rcache_line[2][182].tag_reg.re       = reg2hw.tag_694.re;
  assign rcache_line[2][182].status_reg.status = reg2hw.status_694.q;//status_reg_t'(reg2hw.status_694.q);
  assign rcache_line[2][182].status_reg.qe    = reg2hw.status_694.qe;
  assign rcache_line[2][182].status_reg.re    = reg2hw.status_694.re;


  assign rcache_line[2][183].tag_reg.tag      = reg2hw.tag_695.q;
  assign rcache_line[2][183].tag_reg.qe       = reg2hw.tag_695.qe;
  assign rcache_line[2][183].tag_reg.re       = reg2hw.tag_695.re;
  assign rcache_line[2][183].status_reg.status = reg2hw.status_695.q;//status_reg_t'(reg2hw.status_695.q);
  assign rcache_line[2][183].status_reg.qe    = reg2hw.status_695.qe;
  assign rcache_line[2][183].status_reg.re    = reg2hw.status_695.re;


  assign rcache_line[2][184].tag_reg.tag      = reg2hw.tag_696.q;
  assign rcache_line[2][184].tag_reg.qe       = reg2hw.tag_696.qe;
  assign rcache_line[2][184].tag_reg.re       = reg2hw.tag_696.re;
  assign rcache_line[2][184].status_reg.status = reg2hw.status_696.q;//status_reg_t'(reg2hw.status_696.q);
  assign rcache_line[2][184].status_reg.qe    = reg2hw.status_696.qe;
  assign rcache_line[2][184].status_reg.re    = reg2hw.status_696.re;


  assign rcache_line[2][185].tag_reg.tag      = reg2hw.tag_697.q;
  assign rcache_line[2][185].tag_reg.qe       = reg2hw.tag_697.qe;
  assign rcache_line[2][185].tag_reg.re       = reg2hw.tag_697.re;
  assign rcache_line[2][185].status_reg.status = reg2hw.status_697.q;//status_reg_t'(reg2hw.status_697.q);
  assign rcache_line[2][185].status_reg.qe    = reg2hw.status_697.qe;
  assign rcache_line[2][185].status_reg.re    = reg2hw.status_697.re;


  assign rcache_line[2][186].tag_reg.tag      = reg2hw.tag_698.q;
  assign rcache_line[2][186].tag_reg.qe       = reg2hw.tag_698.qe;
  assign rcache_line[2][186].tag_reg.re       = reg2hw.tag_698.re;
  assign rcache_line[2][186].status_reg.status = reg2hw.status_698.q;//status_reg_t'(reg2hw.status_698.q);
  assign rcache_line[2][186].status_reg.qe    = reg2hw.status_698.qe;
  assign rcache_line[2][186].status_reg.re    = reg2hw.status_698.re;


  assign rcache_line[2][187].tag_reg.tag      = reg2hw.tag_699.q;
  assign rcache_line[2][187].tag_reg.qe       = reg2hw.tag_699.qe;
  assign rcache_line[2][187].tag_reg.re       = reg2hw.tag_699.re;
  assign rcache_line[2][187].status_reg.status = reg2hw.status_699.q;//status_reg_t'(reg2hw.status_699.q);
  assign rcache_line[2][187].status_reg.qe    = reg2hw.status_699.qe;
  assign rcache_line[2][187].status_reg.re    = reg2hw.status_699.re;


  assign rcache_line[2][188].tag_reg.tag      = reg2hw.tag_700.q;
  assign rcache_line[2][188].tag_reg.qe       = reg2hw.tag_700.qe;
  assign rcache_line[2][188].tag_reg.re       = reg2hw.tag_700.re;
  assign rcache_line[2][188].status_reg.status = reg2hw.status_700.q;//status_reg_t'(reg2hw.status_700.q);
  assign rcache_line[2][188].status_reg.qe    = reg2hw.status_700.qe;
  assign rcache_line[2][188].status_reg.re    = reg2hw.status_700.re;


  assign rcache_line[2][189].tag_reg.tag      = reg2hw.tag_701.q;
  assign rcache_line[2][189].tag_reg.qe       = reg2hw.tag_701.qe;
  assign rcache_line[2][189].tag_reg.re       = reg2hw.tag_701.re;
  assign rcache_line[2][189].status_reg.status = reg2hw.status_701.q;//status_reg_t'(reg2hw.status_701.q);
  assign rcache_line[2][189].status_reg.qe    = reg2hw.status_701.qe;
  assign rcache_line[2][189].status_reg.re    = reg2hw.status_701.re;


  assign rcache_line[2][190].tag_reg.tag      = reg2hw.tag_702.q;
  assign rcache_line[2][190].tag_reg.qe       = reg2hw.tag_702.qe;
  assign rcache_line[2][190].tag_reg.re       = reg2hw.tag_702.re;
  assign rcache_line[2][190].status_reg.status = reg2hw.status_702.q;//status_reg_t'(reg2hw.status_702.q);
  assign rcache_line[2][190].status_reg.qe    = reg2hw.status_702.qe;
  assign rcache_line[2][190].status_reg.re    = reg2hw.status_702.re;


  assign rcache_line[2][191].tag_reg.tag      = reg2hw.tag_703.q;
  assign rcache_line[2][191].tag_reg.qe       = reg2hw.tag_703.qe;
  assign rcache_line[2][191].tag_reg.re       = reg2hw.tag_703.re;
  assign rcache_line[2][191].status_reg.status = reg2hw.status_703.q;//status_reg_t'(reg2hw.status_703.q);
  assign rcache_line[2][191].status_reg.qe    = reg2hw.status_703.qe;
  assign rcache_line[2][191].status_reg.re    = reg2hw.status_703.re;


  assign rcache_line[2][192].tag_reg.tag      = reg2hw.tag_704.q;
  assign rcache_line[2][192].tag_reg.qe       = reg2hw.tag_704.qe;
  assign rcache_line[2][192].tag_reg.re       = reg2hw.tag_704.re;
  assign rcache_line[2][192].status_reg.status = reg2hw.status_704.q;//status_reg_t'(reg2hw.status_704.q);
  assign rcache_line[2][192].status_reg.qe    = reg2hw.status_704.qe;
  assign rcache_line[2][192].status_reg.re    = reg2hw.status_704.re;


  assign rcache_line[2][193].tag_reg.tag      = reg2hw.tag_705.q;
  assign rcache_line[2][193].tag_reg.qe       = reg2hw.tag_705.qe;
  assign rcache_line[2][193].tag_reg.re       = reg2hw.tag_705.re;
  assign rcache_line[2][193].status_reg.status = reg2hw.status_705.q;//status_reg_t'(reg2hw.status_705.q);
  assign rcache_line[2][193].status_reg.qe    = reg2hw.status_705.qe;
  assign rcache_line[2][193].status_reg.re    = reg2hw.status_705.re;


  assign rcache_line[2][194].tag_reg.tag      = reg2hw.tag_706.q;
  assign rcache_line[2][194].tag_reg.qe       = reg2hw.tag_706.qe;
  assign rcache_line[2][194].tag_reg.re       = reg2hw.tag_706.re;
  assign rcache_line[2][194].status_reg.status = reg2hw.status_706.q;//status_reg_t'(reg2hw.status_706.q);
  assign rcache_line[2][194].status_reg.qe    = reg2hw.status_706.qe;
  assign rcache_line[2][194].status_reg.re    = reg2hw.status_706.re;


  assign rcache_line[2][195].tag_reg.tag      = reg2hw.tag_707.q;
  assign rcache_line[2][195].tag_reg.qe       = reg2hw.tag_707.qe;
  assign rcache_line[2][195].tag_reg.re       = reg2hw.tag_707.re;
  assign rcache_line[2][195].status_reg.status = reg2hw.status_707.q;//status_reg_t'(reg2hw.status_707.q);
  assign rcache_line[2][195].status_reg.qe    = reg2hw.status_707.qe;
  assign rcache_line[2][195].status_reg.re    = reg2hw.status_707.re;


  assign rcache_line[2][196].tag_reg.tag      = reg2hw.tag_708.q;
  assign rcache_line[2][196].tag_reg.qe       = reg2hw.tag_708.qe;
  assign rcache_line[2][196].tag_reg.re       = reg2hw.tag_708.re;
  assign rcache_line[2][196].status_reg.status = reg2hw.status_708.q;//status_reg_t'(reg2hw.status_708.q);
  assign rcache_line[2][196].status_reg.qe    = reg2hw.status_708.qe;
  assign rcache_line[2][196].status_reg.re    = reg2hw.status_708.re;


  assign rcache_line[2][197].tag_reg.tag      = reg2hw.tag_709.q;
  assign rcache_line[2][197].tag_reg.qe       = reg2hw.tag_709.qe;
  assign rcache_line[2][197].tag_reg.re       = reg2hw.tag_709.re;
  assign rcache_line[2][197].status_reg.status = reg2hw.status_709.q;//status_reg_t'(reg2hw.status_709.q);
  assign rcache_line[2][197].status_reg.qe    = reg2hw.status_709.qe;
  assign rcache_line[2][197].status_reg.re    = reg2hw.status_709.re;


  assign rcache_line[2][198].tag_reg.tag      = reg2hw.tag_710.q;
  assign rcache_line[2][198].tag_reg.qe       = reg2hw.tag_710.qe;
  assign rcache_line[2][198].tag_reg.re       = reg2hw.tag_710.re;
  assign rcache_line[2][198].status_reg.status = reg2hw.status_710.q;//status_reg_t'(reg2hw.status_710.q);
  assign rcache_line[2][198].status_reg.qe    = reg2hw.status_710.qe;
  assign rcache_line[2][198].status_reg.re    = reg2hw.status_710.re;


  assign rcache_line[2][199].tag_reg.tag      = reg2hw.tag_711.q;
  assign rcache_line[2][199].tag_reg.qe       = reg2hw.tag_711.qe;
  assign rcache_line[2][199].tag_reg.re       = reg2hw.tag_711.re;
  assign rcache_line[2][199].status_reg.status = reg2hw.status_711.q;//status_reg_t'(reg2hw.status_711.q);
  assign rcache_line[2][199].status_reg.qe    = reg2hw.status_711.qe;
  assign rcache_line[2][199].status_reg.re    = reg2hw.status_711.re;


  assign rcache_line[2][200].tag_reg.tag      = reg2hw.tag_712.q;
  assign rcache_line[2][200].tag_reg.qe       = reg2hw.tag_712.qe;
  assign rcache_line[2][200].tag_reg.re       = reg2hw.tag_712.re;
  assign rcache_line[2][200].status_reg.status = reg2hw.status_712.q;//status_reg_t'(reg2hw.status_712.q);
  assign rcache_line[2][200].status_reg.qe    = reg2hw.status_712.qe;
  assign rcache_line[2][200].status_reg.re    = reg2hw.status_712.re;


  assign rcache_line[2][201].tag_reg.tag      = reg2hw.tag_713.q;
  assign rcache_line[2][201].tag_reg.qe       = reg2hw.tag_713.qe;
  assign rcache_line[2][201].tag_reg.re       = reg2hw.tag_713.re;
  assign rcache_line[2][201].status_reg.status = reg2hw.status_713.q;//status_reg_t'(reg2hw.status_713.q);
  assign rcache_line[2][201].status_reg.qe    = reg2hw.status_713.qe;
  assign rcache_line[2][201].status_reg.re    = reg2hw.status_713.re;


  assign rcache_line[2][202].tag_reg.tag      = reg2hw.tag_714.q;
  assign rcache_line[2][202].tag_reg.qe       = reg2hw.tag_714.qe;
  assign rcache_line[2][202].tag_reg.re       = reg2hw.tag_714.re;
  assign rcache_line[2][202].status_reg.status = reg2hw.status_714.q;//status_reg_t'(reg2hw.status_714.q);
  assign rcache_line[2][202].status_reg.qe    = reg2hw.status_714.qe;
  assign rcache_line[2][202].status_reg.re    = reg2hw.status_714.re;


  assign rcache_line[2][203].tag_reg.tag      = reg2hw.tag_715.q;
  assign rcache_line[2][203].tag_reg.qe       = reg2hw.tag_715.qe;
  assign rcache_line[2][203].tag_reg.re       = reg2hw.tag_715.re;
  assign rcache_line[2][203].status_reg.status = reg2hw.status_715.q;//status_reg_t'(reg2hw.status_715.q);
  assign rcache_line[2][203].status_reg.qe    = reg2hw.status_715.qe;
  assign rcache_line[2][203].status_reg.re    = reg2hw.status_715.re;


  assign rcache_line[2][204].tag_reg.tag      = reg2hw.tag_716.q;
  assign rcache_line[2][204].tag_reg.qe       = reg2hw.tag_716.qe;
  assign rcache_line[2][204].tag_reg.re       = reg2hw.tag_716.re;
  assign rcache_line[2][204].status_reg.status = reg2hw.status_716.q;//status_reg_t'(reg2hw.status_716.q);
  assign rcache_line[2][204].status_reg.qe    = reg2hw.status_716.qe;
  assign rcache_line[2][204].status_reg.re    = reg2hw.status_716.re;


  assign rcache_line[2][205].tag_reg.tag      = reg2hw.tag_717.q;
  assign rcache_line[2][205].tag_reg.qe       = reg2hw.tag_717.qe;
  assign rcache_line[2][205].tag_reg.re       = reg2hw.tag_717.re;
  assign rcache_line[2][205].status_reg.status = reg2hw.status_717.q;//status_reg_t'(reg2hw.status_717.q);
  assign rcache_line[2][205].status_reg.qe    = reg2hw.status_717.qe;
  assign rcache_line[2][205].status_reg.re    = reg2hw.status_717.re;


  assign rcache_line[2][206].tag_reg.tag      = reg2hw.tag_718.q;
  assign rcache_line[2][206].tag_reg.qe       = reg2hw.tag_718.qe;
  assign rcache_line[2][206].tag_reg.re       = reg2hw.tag_718.re;
  assign rcache_line[2][206].status_reg.status = reg2hw.status_718.q;//status_reg_t'(reg2hw.status_718.q);
  assign rcache_line[2][206].status_reg.qe    = reg2hw.status_718.qe;
  assign rcache_line[2][206].status_reg.re    = reg2hw.status_718.re;


  assign rcache_line[2][207].tag_reg.tag      = reg2hw.tag_719.q;
  assign rcache_line[2][207].tag_reg.qe       = reg2hw.tag_719.qe;
  assign rcache_line[2][207].tag_reg.re       = reg2hw.tag_719.re;
  assign rcache_line[2][207].status_reg.status = reg2hw.status_719.q;//status_reg_t'(reg2hw.status_719.q);
  assign rcache_line[2][207].status_reg.qe    = reg2hw.status_719.qe;
  assign rcache_line[2][207].status_reg.re    = reg2hw.status_719.re;


  assign rcache_line[2][208].tag_reg.tag      = reg2hw.tag_720.q;
  assign rcache_line[2][208].tag_reg.qe       = reg2hw.tag_720.qe;
  assign rcache_line[2][208].tag_reg.re       = reg2hw.tag_720.re;
  assign rcache_line[2][208].status_reg.status = reg2hw.status_720.q;//status_reg_t'(reg2hw.status_720.q);
  assign rcache_line[2][208].status_reg.qe    = reg2hw.status_720.qe;
  assign rcache_line[2][208].status_reg.re    = reg2hw.status_720.re;


  assign rcache_line[2][209].tag_reg.tag      = reg2hw.tag_721.q;
  assign rcache_line[2][209].tag_reg.qe       = reg2hw.tag_721.qe;
  assign rcache_line[2][209].tag_reg.re       = reg2hw.tag_721.re;
  assign rcache_line[2][209].status_reg.status = reg2hw.status_721.q;//status_reg_t'(reg2hw.status_721.q);
  assign rcache_line[2][209].status_reg.qe    = reg2hw.status_721.qe;
  assign rcache_line[2][209].status_reg.re    = reg2hw.status_721.re;


  assign rcache_line[2][210].tag_reg.tag      = reg2hw.tag_722.q;
  assign rcache_line[2][210].tag_reg.qe       = reg2hw.tag_722.qe;
  assign rcache_line[2][210].tag_reg.re       = reg2hw.tag_722.re;
  assign rcache_line[2][210].status_reg.status = reg2hw.status_722.q;//status_reg_t'(reg2hw.status_722.q);
  assign rcache_line[2][210].status_reg.qe    = reg2hw.status_722.qe;
  assign rcache_line[2][210].status_reg.re    = reg2hw.status_722.re;


  assign rcache_line[2][211].tag_reg.tag      = reg2hw.tag_723.q;
  assign rcache_line[2][211].tag_reg.qe       = reg2hw.tag_723.qe;
  assign rcache_line[2][211].tag_reg.re       = reg2hw.tag_723.re;
  assign rcache_line[2][211].status_reg.status = reg2hw.status_723.q;//status_reg_t'(reg2hw.status_723.q);
  assign rcache_line[2][211].status_reg.qe    = reg2hw.status_723.qe;
  assign rcache_line[2][211].status_reg.re    = reg2hw.status_723.re;


  assign rcache_line[2][212].tag_reg.tag      = reg2hw.tag_724.q;
  assign rcache_line[2][212].tag_reg.qe       = reg2hw.tag_724.qe;
  assign rcache_line[2][212].tag_reg.re       = reg2hw.tag_724.re;
  assign rcache_line[2][212].status_reg.status = reg2hw.status_724.q;//status_reg_t'(reg2hw.status_724.q);
  assign rcache_line[2][212].status_reg.qe    = reg2hw.status_724.qe;
  assign rcache_line[2][212].status_reg.re    = reg2hw.status_724.re;


  assign rcache_line[2][213].tag_reg.tag      = reg2hw.tag_725.q;
  assign rcache_line[2][213].tag_reg.qe       = reg2hw.tag_725.qe;
  assign rcache_line[2][213].tag_reg.re       = reg2hw.tag_725.re;
  assign rcache_line[2][213].status_reg.status = reg2hw.status_725.q;//status_reg_t'(reg2hw.status_725.q);
  assign rcache_line[2][213].status_reg.qe    = reg2hw.status_725.qe;
  assign rcache_line[2][213].status_reg.re    = reg2hw.status_725.re;


  assign rcache_line[2][214].tag_reg.tag      = reg2hw.tag_726.q;
  assign rcache_line[2][214].tag_reg.qe       = reg2hw.tag_726.qe;
  assign rcache_line[2][214].tag_reg.re       = reg2hw.tag_726.re;
  assign rcache_line[2][214].status_reg.status = reg2hw.status_726.q;//status_reg_t'(reg2hw.status_726.q);
  assign rcache_line[2][214].status_reg.qe    = reg2hw.status_726.qe;
  assign rcache_line[2][214].status_reg.re    = reg2hw.status_726.re;


  assign rcache_line[2][215].tag_reg.tag      = reg2hw.tag_727.q;
  assign rcache_line[2][215].tag_reg.qe       = reg2hw.tag_727.qe;
  assign rcache_line[2][215].tag_reg.re       = reg2hw.tag_727.re;
  assign rcache_line[2][215].status_reg.status = reg2hw.status_727.q;//status_reg_t'(reg2hw.status_727.q);
  assign rcache_line[2][215].status_reg.qe    = reg2hw.status_727.qe;
  assign rcache_line[2][215].status_reg.re    = reg2hw.status_727.re;


  assign rcache_line[2][216].tag_reg.tag      = reg2hw.tag_728.q;
  assign rcache_line[2][216].tag_reg.qe       = reg2hw.tag_728.qe;
  assign rcache_line[2][216].tag_reg.re       = reg2hw.tag_728.re;
  assign rcache_line[2][216].status_reg.status = reg2hw.status_728.q;//status_reg_t'(reg2hw.status_728.q);
  assign rcache_line[2][216].status_reg.qe    = reg2hw.status_728.qe;
  assign rcache_line[2][216].status_reg.re    = reg2hw.status_728.re;


  assign rcache_line[2][217].tag_reg.tag      = reg2hw.tag_729.q;
  assign rcache_line[2][217].tag_reg.qe       = reg2hw.tag_729.qe;
  assign rcache_line[2][217].tag_reg.re       = reg2hw.tag_729.re;
  assign rcache_line[2][217].status_reg.status = reg2hw.status_729.q;//status_reg_t'(reg2hw.status_729.q);
  assign rcache_line[2][217].status_reg.qe    = reg2hw.status_729.qe;
  assign rcache_line[2][217].status_reg.re    = reg2hw.status_729.re;


  assign rcache_line[2][218].tag_reg.tag      = reg2hw.tag_730.q;
  assign rcache_line[2][218].tag_reg.qe       = reg2hw.tag_730.qe;
  assign rcache_line[2][218].tag_reg.re       = reg2hw.tag_730.re;
  assign rcache_line[2][218].status_reg.status = reg2hw.status_730.q;//status_reg_t'(reg2hw.status_730.q);
  assign rcache_line[2][218].status_reg.qe    = reg2hw.status_730.qe;
  assign rcache_line[2][218].status_reg.re    = reg2hw.status_730.re;


  assign rcache_line[2][219].tag_reg.tag      = reg2hw.tag_731.q;
  assign rcache_line[2][219].tag_reg.qe       = reg2hw.tag_731.qe;
  assign rcache_line[2][219].tag_reg.re       = reg2hw.tag_731.re;
  assign rcache_line[2][219].status_reg.status = reg2hw.status_731.q;//status_reg_t'(reg2hw.status_731.q);
  assign rcache_line[2][219].status_reg.qe    = reg2hw.status_731.qe;
  assign rcache_line[2][219].status_reg.re    = reg2hw.status_731.re;


  assign rcache_line[2][220].tag_reg.tag      = reg2hw.tag_732.q;
  assign rcache_line[2][220].tag_reg.qe       = reg2hw.tag_732.qe;
  assign rcache_line[2][220].tag_reg.re       = reg2hw.tag_732.re;
  assign rcache_line[2][220].status_reg.status = reg2hw.status_732.q;//status_reg_t'(reg2hw.status_732.q);
  assign rcache_line[2][220].status_reg.qe    = reg2hw.status_732.qe;
  assign rcache_line[2][220].status_reg.re    = reg2hw.status_732.re;


  assign rcache_line[2][221].tag_reg.tag      = reg2hw.tag_733.q;
  assign rcache_line[2][221].tag_reg.qe       = reg2hw.tag_733.qe;
  assign rcache_line[2][221].tag_reg.re       = reg2hw.tag_733.re;
  assign rcache_line[2][221].status_reg.status = reg2hw.status_733.q;//status_reg_t'(reg2hw.status_733.q);
  assign rcache_line[2][221].status_reg.qe    = reg2hw.status_733.qe;
  assign rcache_line[2][221].status_reg.re    = reg2hw.status_733.re;


  assign rcache_line[2][222].tag_reg.tag      = reg2hw.tag_734.q;
  assign rcache_line[2][222].tag_reg.qe       = reg2hw.tag_734.qe;
  assign rcache_line[2][222].tag_reg.re       = reg2hw.tag_734.re;
  assign rcache_line[2][222].status_reg.status = reg2hw.status_734.q;//status_reg_t'(reg2hw.status_734.q);
  assign rcache_line[2][222].status_reg.qe    = reg2hw.status_734.qe;
  assign rcache_line[2][222].status_reg.re    = reg2hw.status_734.re;


  assign rcache_line[2][223].tag_reg.tag      = reg2hw.tag_735.q;
  assign rcache_line[2][223].tag_reg.qe       = reg2hw.tag_735.qe;
  assign rcache_line[2][223].tag_reg.re       = reg2hw.tag_735.re;
  assign rcache_line[2][223].status_reg.status = reg2hw.status_735.q;//status_reg_t'(reg2hw.status_735.q);
  assign rcache_line[2][223].status_reg.qe    = reg2hw.status_735.qe;
  assign rcache_line[2][223].status_reg.re    = reg2hw.status_735.re;


  assign rcache_line[2][224].tag_reg.tag      = reg2hw.tag_736.q;
  assign rcache_line[2][224].tag_reg.qe       = reg2hw.tag_736.qe;
  assign rcache_line[2][224].tag_reg.re       = reg2hw.tag_736.re;
  assign rcache_line[2][224].status_reg.status = reg2hw.status_736.q;//status_reg_t'(reg2hw.status_736.q);
  assign rcache_line[2][224].status_reg.qe    = reg2hw.status_736.qe;
  assign rcache_line[2][224].status_reg.re    = reg2hw.status_736.re;


  assign rcache_line[2][225].tag_reg.tag      = reg2hw.tag_737.q;
  assign rcache_line[2][225].tag_reg.qe       = reg2hw.tag_737.qe;
  assign rcache_line[2][225].tag_reg.re       = reg2hw.tag_737.re;
  assign rcache_line[2][225].status_reg.status = reg2hw.status_737.q;//status_reg_t'(reg2hw.status_737.q);
  assign rcache_line[2][225].status_reg.qe    = reg2hw.status_737.qe;
  assign rcache_line[2][225].status_reg.re    = reg2hw.status_737.re;


  assign rcache_line[2][226].tag_reg.tag      = reg2hw.tag_738.q;
  assign rcache_line[2][226].tag_reg.qe       = reg2hw.tag_738.qe;
  assign rcache_line[2][226].tag_reg.re       = reg2hw.tag_738.re;
  assign rcache_line[2][226].status_reg.status = reg2hw.status_738.q;//status_reg_t'(reg2hw.status_738.q);
  assign rcache_line[2][226].status_reg.qe    = reg2hw.status_738.qe;
  assign rcache_line[2][226].status_reg.re    = reg2hw.status_738.re;


  assign rcache_line[2][227].tag_reg.tag      = reg2hw.tag_739.q;
  assign rcache_line[2][227].tag_reg.qe       = reg2hw.tag_739.qe;
  assign rcache_line[2][227].tag_reg.re       = reg2hw.tag_739.re;
  assign rcache_line[2][227].status_reg.status = reg2hw.status_739.q;//status_reg_t'(reg2hw.status_739.q);
  assign rcache_line[2][227].status_reg.qe    = reg2hw.status_739.qe;
  assign rcache_line[2][227].status_reg.re    = reg2hw.status_739.re;


  assign rcache_line[2][228].tag_reg.tag      = reg2hw.tag_740.q;
  assign rcache_line[2][228].tag_reg.qe       = reg2hw.tag_740.qe;
  assign rcache_line[2][228].tag_reg.re       = reg2hw.tag_740.re;
  assign rcache_line[2][228].status_reg.status = reg2hw.status_740.q;//status_reg_t'(reg2hw.status_740.q);
  assign rcache_line[2][228].status_reg.qe    = reg2hw.status_740.qe;
  assign rcache_line[2][228].status_reg.re    = reg2hw.status_740.re;


  assign rcache_line[2][229].tag_reg.tag      = reg2hw.tag_741.q;
  assign rcache_line[2][229].tag_reg.qe       = reg2hw.tag_741.qe;
  assign rcache_line[2][229].tag_reg.re       = reg2hw.tag_741.re;
  assign rcache_line[2][229].status_reg.status = reg2hw.status_741.q;//status_reg_t'(reg2hw.status_741.q);
  assign rcache_line[2][229].status_reg.qe    = reg2hw.status_741.qe;
  assign rcache_line[2][229].status_reg.re    = reg2hw.status_741.re;


  assign rcache_line[2][230].tag_reg.tag      = reg2hw.tag_742.q;
  assign rcache_line[2][230].tag_reg.qe       = reg2hw.tag_742.qe;
  assign rcache_line[2][230].tag_reg.re       = reg2hw.tag_742.re;
  assign rcache_line[2][230].status_reg.status = reg2hw.status_742.q;//status_reg_t'(reg2hw.status_742.q);
  assign rcache_line[2][230].status_reg.qe    = reg2hw.status_742.qe;
  assign rcache_line[2][230].status_reg.re    = reg2hw.status_742.re;


  assign rcache_line[2][231].tag_reg.tag      = reg2hw.tag_743.q;
  assign rcache_line[2][231].tag_reg.qe       = reg2hw.tag_743.qe;
  assign rcache_line[2][231].tag_reg.re       = reg2hw.tag_743.re;
  assign rcache_line[2][231].status_reg.status = reg2hw.status_743.q;//status_reg_t'(reg2hw.status_743.q);
  assign rcache_line[2][231].status_reg.qe    = reg2hw.status_743.qe;
  assign rcache_line[2][231].status_reg.re    = reg2hw.status_743.re;


  assign rcache_line[2][232].tag_reg.tag      = reg2hw.tag_744.q;
  assign rcache_line[2][232].tag_reg.qe       = reg2hw.tag_744.qe;
  assign rcache_line[2][232].tag_reg.re       = reg2hw.tag_744.re;
  assign rcache_line[2][232].status_reg.status = reg2hw.status_744.q;//status_reg_t'(reg2hw.status_744.q);
  assign rcache_line[2][232].status_reg.qe    = reg2hw.status_744.qe;
  assign rcache_line[2][232].status_reg.re    = reg2hw.status_744.re;


  assign rcache_line[2][233].tag_reg.tag      = reg2hw.tag_745.q;
  assign rcache_line[2][233].tag_reg.qe       = reg2hw.tag_745.qe;
  assign rcache_line[2][233].tag_reg.re       = reg2hw.tag_745.re;
  assign rcache_line[2][233].status_reg.status = reg2hw.status_745.q;//status_reg_t'(reg2hw.status_745.q);
  assign rcache_line[2][233].status_reg.qe    = reg2hw.status_745.qe;
  assign rcache_line[2][233].status_reg.re    = reg2hw.status_745.re;


  assign rcache_line[2][234].tag_reg.tag      = reg2hw.tag_746.q;
  assign rcache_line[2][234].tag_reg.qe       = reg2hw.tag_746.qe;
  assign rcache_line[2][234].tag_reg.re       = reg2hw.tag_746.re;
  assign rcache_line[2][234].status_reg.status = reg2hw.status_746.q;//status_reg_t'(reg2hw.status_746.q);
  assign rcache_line[2][234].status_reg.qe    = reg2hw.status_746.qe;
  assign rcache_line[2][234].status_reg.re    = reg2hw.status_746.re;


  assign rcache_line[2][235].tag_reg.tag      = reg2hw.tag_747.q;
  assign rcache_line[2][235].tag_reg.qe       = reg2hw.tag_747.qe;
  assign rcache_line[2][235].tag_reg.re       = reg2hw.tag_747.re;
  assign rcache_line[2][235].status_reg.status = reg2hw.status_747.q;//status_reg_t'(reg2hw.status_747.q);
  assign rcache_line[2][235].status_reg.qe    = reg2hw.status_747.qe;
  assign rcache_line[2][235].status_reg.re    = reg2hw.status_747.re;


  assign rcache_line[2][236].tag_reg.tag      = reg2hw.tag_748.q;
  assign rcache_line[2][236].tag_reg.qe       = reg2hw.tag_748.qe;
  assign rcache_line[2][236].tag_reg.re       = reg2hw.tag_748.re;
  assign rcache_line[2][236].status_reg.status = reg2hw.status_748.q;//status_reg_t'(reg2hw.status_748.q);
  assign rcache_line[2][236].status_reg.qe    = reg2hw.status_748.qe;
  assign rcache_line[2][236].status_reg.re    = reg2hw.status_748.re;


  assign rcache_line[2][237].tag_reg.tag      = reg2hw.tag_749.q;
  assign rcache_line[2][237].tag_reg.qe       = reg2hw.tag_749.qe;
  assign rcache_line[2][237].tag_reg.re       = reg2hw.tag_749.re;
  assign rcache_line[2][237].status_reg.status = reg2hw.status_749.q;//status_reg_t'(reg2hw.status_749.q);
  assign rcache_line[2][237].status_reg.qe    = reg2hw.status_749.qe;
  assign rcache_line[2][237].status_reg.re    = reg2hw.status_749.re;


  assign rcache_line[2][238].tag_reg.tag      = reg2hw.tag_750.q;
  assign rcache_line[2][238].tag_reg.qe       = reg2hw.tag_750.qe;
  assign rcache_line[2][238].tag_reg.re       = reg2hw.tag_750.re;
  assign rcache_line[2][238].status_reg.status = reg2hw.status_750.q;//status_reg_t'(reg2hw.status_750.q);
  assign rcache_line[2][238].status_reg.qe    = reg2hw.status_750.qe;
  assign rcache_line[2][238].status_reg.re    = reg2hw.status_750.re;


  assign rcache_line[2][239].tag_reg.tag      = reg2hw.tag_751.q;
  assign rcache_line[2][239].tag_reg.qe       = reg2hw.tag_751.qe;
  assign rcache_line[2][239].tag_reg.re       = reg2hw.tag_751.re;
  assign rcache_line[2][239].status_reg.status = reg2hw.status_751.q;//status_reg_t'(reg2hw.status_751.q);
  assign rcache_line[2][239].status_reg.qe    = reg2hw.status_751.qe;
  assign rcache_line[2][239].status_reg.re    = reg2hw.status_751.re;


  assign rcache_line[2][240].tag_reg.tag      = reg2hw.tag_752.q;
  assign rcache_line[2][240].tag_reg.qe       = reg2hw.tag_752.qe;
  assign rcache_line[2][240].tag_reg.re       = reg2hw.tag_752.re;
  assign rcache_line[2][240].status_reg.status = reg2hw.status_752.q;//status_reg_t'(reg2hw.status_752.q);
  assign rcache_line[2][240].status_reg.qe    = reg2hw.status_752.qe;
  assign rcache_line[2][240].status_reg.re    = reg2hw.status_752.re;


  assign rcache_line[2][241].tag_reg.tag      = reg2hw.tag_753.q;
  assign rcache_line[2][241].tag_reg.qe       = reg2hw.tag_753.qe;
  assign rcache_line[2][241].tag_reg.re       = reg2hw.tag_753.re;
  assign rcache_line[2][241].status_reg.status = reg2hw.status_753.q;//status_reg_t'(reg2hw.status_753.q);
  assign rcache_line[2][241].status_reg.qe    = reg2hw.status_753.qe;
  assign rcache_line[2][241].status_reg.re    = reg2hw.status_753.re;


  assign rcache_line[2][242].tag_reg.tag      = reg2hw.tag_754.q;
  assign rcache_line[2][242].tag_reg.qe       = reg2hw.tag_754.qe;
  assign rcache_line[2][242].tag_reg.re       = reg2hw.tag_754.re;
  assign rcache_line[2][242].status_reg.status = reg2hw.status_754.q;//status_reg_t'(reg2hw.status_754.q);
  assign rcache_line[2][242].status_reg.qe    = reg2hw.status_754.qe;
  assign rcache_line[2][242].status_reg.re    = reg2hw.status_754.re;


  assign rcache_line[2][243].tag_reg.tag      = reg2hw.tag_755.q;
  assign rcache_line[2][243].tag_reg.qe       = reg2hw.tag_755.qe;
  assign rcache_line[2][243].tag_reg.re       = reg2hw.tag_755.re;
  assign rcache_line[2][243].status_reg.status = reg2hw.status_755.q;//status_reg_t'(reg2hw.status_755.q);
  assign rcache_line[2][243].status_reg.qe    = reg2hw.status_755.qe;
  assign rcache_line[2][243].status_reg.re    = reg2hw.status_755.re;


  assign rcache_line[2][244].tag_reg.tag      = reg2hw.tag_756.q;
  assign rcache_line[2][244].tag_reg.qe       = reg2hw.tag_756.qe;
  assign rcache_line[2][244].tag_reg.re       = reg2hw.tag_756.re;
  assign rcache_line[2][244].status_reg.status = reg2hw.status_756.q;//status_reg_t'(reg2hw.status_756.q);
  assign rcache_line[2][244].status_reg.qe    = reg2hw.status_756.qe;
  assign rcache_line[2][244].status_reg.re    = reg2hw.status_756.re;


  assign rcache_line[2][245].tag_reg.tag      = reg2hw.tag_757.q;
  assign rcache_line[2][245].tag_reg.qe       = reg2hw.tag_757.qe;
  assign rcache_line[2][245].tag_reg.re       = reg2hw.tag_757.re;
  assign rcache_line[2][245].status_reg.status = reg2hw.status_757.q;//status_reg_t'(reg2hw.status_757.q);
  assign rcache_line[2][245].status_reg.qe    = reg2hw.status_757.qe;
  assign rcache_line[2][245].status_reg.re    = reg2hw.status_757.re;


  assign rcache_line[2][246].tag_reg.tag      = reg2hw.tag_758.q;
  assign rcache_line[2][246].tag_reg.qe       = reg2hw.tag_758.qe;
  assign rcache_line[2][246].tag_reg.re       = reg2hw.tag_758.re;
  assign rcache_line[2][246].status_reg.status = reg2hw.status_758.q;//status_reg_t'(reg2hw.status_758.q);
  assign rcache_line[2][246].status_reg.qe    = reg2hw.status_758.qe;
  assign rcache_line[2][246].status_reg.re    = reg2hw.status_758.re;


  assign rcache_line[2][247].tag_reg.tag      = reg2hw.tag_759.q;
  assign rcache_line[2][247].tag_reg.qe       = reg2hw.tag_759.qe;
  assign rcache_line[2][247].tag_reg.re       = reg2hw.tag_759.re;
  assign rcache_line[2][247].status_reg.status = reg2hw.status_759.q;//status_reg_t'(reg2hw.status_759.q);
  assign rcache_line[2][247].status_reg.qe    = reg2hw.status_759.qe;
  assign rcache_line[2][247].status_reg.re    = reg2hw.status_759.re;


  assign rcache_line[2][248].tag_reg.tag      = reg2hw.tag_760.q;
  assign rcache_line[2][248].tag_reg.qe       = reg2hw.tag_760.qe;
  assign rcache_line[2][248].tag_reg.re       = reg2hw.tag_760.re;
  assign rcache_line[2][248].status_reg.status = reg2hw.status_760.q;//status_reg_t'(reg2hw.status_760.q);
  assign rcache_line[2][248].status_reg.qe    = reg2hw.status_760.qe;
  assign rcache_line[2][248].status_reg.re    = reg2hw.status_760.re;


  assign rcache_line[2][249].tag_reg.tag      = reg2hw.tag_761.q;
  assign rcache_line[2][249].tag_reg.qe       = reg2hw.tag_761.qe;
  assign rcache_line[2][249].tag_reg.re       = reg2hw.tag_761.re;
  assign rcache_line[2][249].status_reg.status = reg2hw.status_761.q;//status_reg_t'(reg2hw.status_761.q);
  assign rcache_line[2][249].status_reg.qe    = reg2hw.status_761.qe;
  assign rcache_line[2][249].status_reg.re    = reg2hw.status_761.re;


  assign rcache_line[2][250].tag_reg.tag      = reg2hw.tag_762.q;
  assign rcache_line[2][250].tag_reg.qe       = reg2hw.tag_762.qe;
  assign rcache_line[2][250].tag_reg.re       = reg2hw.tag_762.re;
  assign rcache_line[2][250].status_reg.status = reg2hw.status_762.q;//status_reg_t'(reg2hw.status_762.q);
  assign rcache_line[2][250].status_reg.qe    = reg2hw.status_762.qe;
  assign rcache_line[2][250].status_reg.re    = reg2hw.status_762.re;


  assign rcache_line[2][251].tag_reg.tag      = reg2hw.tag_763.q;
  assign rcache_line[2][251].tag_reg.qe       = reg2hw.tag_763.qe;
  assign rcache_line[2][251].tag_reg.re       = reg2hw.tag_763.re;
  assign rcache_line[2][251].status_reg.status = reg2hw.status_763.q;//status_reg_t'(reg2hw.status_763.q);
  assign rcache_line[2][251].status_reg.qe    = reg2hw.status_763.qe;
  assign rcache_line[2][251].status_reg.re    = reg2hw.status_763.re;


  assign rcache_line[2][252].tag_reg.tag      = reg2hw.tag_764.q;
  assign rcache_line[2][252].tag_reg.qe       = reg2hw.tag_764.qe;
  assign rcache_line[2][252].tag_reg.re       = reg2hw.tag_764.re;
  assign rcache_line[2][252].status_reg.status = reg2hw.status_764.q;//status_reg_t'(reg2hw.status_764.q);
  assign rcache_line[2][252].status_reg.qe    = reg2hw.status_764.qe;
  assign rcache_line[2][252].status_reg.re    = reg2hw.status_764.re;


  assign rcache_line[2][253].tag_reg.tag      = reg2hw.tag_765.q;
  assign rcache_line[2][253].tag_reg.qe       = reg2hw.tag_765.qe;
  assign rcache_line[2][253].tag_reg.re       = reg2hw.tag_765.re;
  assign rcache_line[2][253].status_reg.status = reg2hw.status_765.q;//status_reg_t'(reg2hw.status_765.q);
  assign rcache_line[2][253].status_reg.qe    = reg2hw.status_765.qe;
  assign rcache_line[2][253].status_reg.re    = reg2hw.status_765.re;


  assign rcache_line[2][254].tag_reg.tag      = reg2hw.tag_766.q;
  assign rcache_line[2][254].tag_reg.qe       = reg2hw.tag_766.qe;
  assign rcache_line[2][254].tag_reg.re       = reg2hw.tag_766.re;
  assign rcache_line[2][254].status_reg.status = reg2hw.status_766.q;//status_reg_t'(reg2hw.status_766.q);
  assign rcache_line[2][254].status_reg.qe    = reg2hw.status_766.qe;
  assign rcache_line[2][254].status_reg.re    = reg2hw.status_766.re;


  assign rcache_line[2][255].tag_reg.tag      = reg2hw.tag_767.q;
  assign rcache_line[2][255].tag_reg.qe       = reg2hw.tag_767.qe;
  assign rcache_line[2][255].tag_reg.re       = reg2hw.tag_767.re;
  assign rcache_line[2][255].status_reg.status = reg2hw.status_767.q;//status_reg_t'(reg2hw.status_767.q);
  assign rcache_line[2][255].status_reg.qe    = reg2hw.status_767.qe;
  assign rcache_line[2][255].status_reg.re    = reg2hw.status_767.re;


  assign rcache_line[3][0].tag_reg.tag      = reg2hw.tag_768.q;
  assign rcache_line[3][0].tag_reg.qe       = reg2hw.tag_768.qe;
  assign rcache_line[3][0].tag_reg.re       = reg2hw.tag_768.re;
  assign rcache_line[3][0].status_reg.status = reg2hw.status_768.q;//status_reg_t'(reg2hw.status_768.q);
  assign rcache_line[3][0].status_reg.qe    = reg2hw.status_768.qe;
  assign rcache_line[3][0].status_reg.re    = reg2hw.status_768.re;


  assign rcache_line[3][1].tag_reg.tag      = reg2hw.tag_769.q;
  assign rcache_line[3][1].tag_reg.qe       = reg2hw.tag_769.qe;
  assign rcache_line[3][1].tag_reg.re       = reg2hw.tag_769.re;
  assign rcache_line[3][1].status_reg.status = reg2hw.status_769.q;//status_reg_t'(reg2hw.status_769.q);
  assign rcache_line[3][1].status_reg.qe    = reg2hw.status_769.qe;
  assign rcache_line[3][1].status_reg.re    = reg2hw.status_769.re;


  assign rcache_line[3][2].tag_reg.tag      = reg2hw.tag_770.q;
  assign rcache_line[3][2].tag_reg.qe       = reg2hw.tag_770.qe;
  assign rcache_line[3][2].tag_reg.re       = reg2hw.tag_770.re;
  assign rcache_line[3][2].status_reg.status = reg2hw.status_770.q;//status_reg_t'(reg2hw.status_770.q);
  assign rcache_line[3][2].status_reg.qe    = reg2hw.status_770.qe;
  assign rcache_line[3][2].status_reg.re    = reg2hw.status_770.re;


  assign rcache_line[3][3].tag_reg.tag      = reg2hw.tag_771.q;
  assign rcache_line[3][3].tag_reg.qe       = reg2hw.tag_771.qe;
  assign rcache_line[3][3].tag_reg.re       = reg2hw.tag_771.re;
  assign rcache_line[3][3].status_reg.status = reg2hw.status_771.q;//status_reg_t'(reg2hw.status_771.q);
  assign rcache_line[3][3].status_reg.qe    = reg2hw.status_771.qe;
  assign rcache_line[3][3].status_reg.re    = reg2hw.status_771.re;


  assign rcache_line[3][4].tag_reg.tag      = reg2hw.tag_772.q;
  assign rcache_line[3][4].tag_reg.qe       = reg2hw.tag_772.qe;
  assign rcache_line[3][4].tag_reg.re       = reg2hw.tag_772.re;
  assign rcache_line[3][4].status_reg.status = reg2hw.status_772.q;//status_reg_t'(reg2hw.status_772.q);
  assign rcache_line[3][4].status_reg.qe    = reg2hw.status_772.qe;
  assign rcache_line[3][4].status_reg.re    = reg2hw.status_772.re;


  assign rcache_line[3][5].tag_reg.tag      = reg2hw.tag_773.q;
  assign rcache_line[3][5].tag_reg.qe       = reg2hw.tag_773.qe;
  assign rcache_line[3][5].tag_reg.re       = reg2hw.tag_773.re;
  assign rcache_line[3][5].status_reg.status = reg2hw.status_773.q;//status_reg_t'(reg2hw.status_773.q);
  assign rcache_line[3][5].status_reg.qe    = reg2hw.status_773.qe;
  assign rcache_line[3][5].status_reg.re    = reg2hw.status_773.re;


  assign rcache_line[3][6].tag_reg.tag      = reg2hw.tag_774.q;
  assign rcache_line[3][6].tag_reg.qe       = reg2hw.tag_774.qe;
  assign rcache_line[3][6].tag_reg.re       = reg2hw.tag_774.re;
  assign rcache_line[3][6].status_reg.status = reg2hw.status_774.q;//status_reg_t'(reg2hw.status_774.q);
  assign rcache_line[3][6].status_reg.qe    = reg2hw.status_774.qe;
  assign rcache_line[3][6].status_reg.re    = reg2hw.status_774.re;


  assign rcache_line[3][7].tag_reg.tag      = reg2hw.tag_775.q;
  assign rcache_line[3][7].tag_reg.qe       = reg2hw.tag_775.qe;
  assign rcache_line[3][7].tag_reg.re       = reg2hw.tag_775.re;
  assign rcache_line[3][7].status_reg.status = reg2hw.status_775.q;//status_reg_t'(reg2hw.status_775.q);
  assign rcache_line[3][7].status_reg.qe    = reg2hw.status_775.qe;
  assign rcache_line[3][7].status_reg.re    = reg2hw.status_775.re;


  assign rcache_line[3][8].tag_reg.tag      = reg2hw.tag_776.q;
  assign rcache_line[3][8].tag_reg.qe       = reg2hw.tag_776.qe;
  assign rcache_line[3][8].tag_reg.re       = reg2hw.tag_776.re;
  assign rcache_line[3][8].status_reg.status = reg2hw.status_776.q;//status_reg_t'(reg2hw.status_776.q);
  assign rcache_line[3][8].status_reg.qe    = reg2hw.status_776.qe;
  assign rcache_line[3][8].status_reg.re    = reg2hw.status_776.re;


  assign rcache_line[3][9].tag_reg.tag      = reg2hw.tag_777.q;
  assign rcache_line[3][9].tag_reg.qe       = reg2hw.tag_777.qe;
  assign rcache_line[3][9].tag_reg.re       = reg2hw.tag_777.re;
  assign rcache_line[3][9].status_reg.status = reg2hw.status_777.q;//status_reg_t'(reg2hw.status_777.q);
  assign rcache_line[3][9].status_reg.qe    = reg2hw.status_777.qe;
  assign rcache_line[3][9].status_reg.re    = reg2hw.status_777.re;


  assign rcache_line[3][10].tag_reg.tag      = reg2hw.tag_778.q;
  assign rcache_line[3][10].tag_reg.qe       = reg2hw.tag_778.qe;
  assign rcache_line[3][10].tag_reg.re       = reg2hw.tag_778.re;
  assign rcache_line[3][10].status_reg.status = reg2hw.status_778.q;//status_reg_t'(reg2hw.status_778.q);
  assign rcache_line[3][10].status_reg.qe    = reg2hw.status_778.qe;
  assign rcache_line[3][10].status_reg.re    = reg2hw.status_778.re;


  assign rcache_line[3][11].tag_reg.tag      = reg2hw.tag_779.q;
  assign rcache_line[3][11].tag_reg.qe       = reg2hw.tag_779.qe;
  assign rcache_line[3][11].tag_reg.re       = reg2hw.tag_779.re;
  assign rcache_line[3][11].status_reg.status = reg2hw.status_779.q;//status_reg_t'(reg2hw.status_779.q);
  assign rcache_line[3][11].status_reg.qe    = reg2hw.status_779.qe;
  assign rcache_line[3][11].status_reg.re    = reg2hw.status_779.re;


  assign rcache_line[3][12].tag_reg.tag      = reg2hw.tag_780.q;
  assign rcache_line[3][12].tag_reg.qe       = reg2hw.tag_780.qe;
  assign rcache_line[3][12].tag_reg.re       = reg2hw.tag_780.re;
  assign rcache_line[3][12].status_reg.status = reg2hw.status_780.q;//status_reg_t'(reg2hw.status_780.q);
  assign rcache_line[3][12].status_reg.qe    = reg2hw.status_780.qe;
  assign rcache_line[3][12].status_reg.re    = reg2hw.status_780.re;


  assign rcache_line[3][13].tag_reg.tag      = reg2hw.tag_781.q;
  assign rcache_line[3][13].tag_reg.qe       = reg2hw.tag_781.qe;
  assign rcache_line[3][13].tag_reg.re       = reg2hw.tag_781.re;
  assign rcache_line[3][13].status_reg.status = reg2hw.status_781.q;//status_reg_t'(reg2hw.status_781.q);
  assign rcache_line[3][13].status_reg.qe    = reg2hw.status_781.qe;
  assign rcache_line[3][13].status_reg.re    = reg2hw.status_781.re;


  assign rcache_line[3][14].tag_reg.tag      = reg2hw.tag_782.q;
  assign rcache_line[3][14].tag_reg.qe       = reg2hw.tag_782.qe;
  assign rcache_line[3][14].tag_reg.re       = reg2hw.tag_782.re;
  assign rcache_line[3][14].status_reg.status = reg2hw.status_782.q;//status_reg_t'(reg2hw.status_782.q);
  assign rcache_line[3][14].status_reg.qe    = reg2hw.status_782.qe;
  assign rcache_line[3][14].status_reg.re    = reg2hw.status_782.re;


  assign rcache_line[3][15].tag_reg.tag      = reg2hw.tag_783.q;
  assign rcache_line[3][15].tag_reg.qe       = reg2hw.tag_783.qe;
  assign rcache_line[3][15].tag_reg.re       = reg2hw.tag_783.re;
  assign rcache_line[3][15].status_reg.status = reg2hw.status_783.q;//status_reg_t'(reg2hw.status_783.q);
  assign rcache_line[3][15].status_reg.qe    = reg2hw.status_783.qe;
  assign rcache_line[3][15].status_reg.re    = reg2hw.status_783.re;


  assign rcache_line[3][16].tag_reg.tag      = reg2hw.tag_784.q;
  assign rcache_line[3][16].tag_reg.qe       = reg2hw.tag_784.qe;
  assign rcache_line[3][16].tag_reg.re       = reg2hw.tag_784.re;
  assign rcache_line[3][16].status_reg.status = reg2hw.status_784.q;//status_reg_t'(reg2hw.status_784.q);
  assign rcache_line[3][16].status_reg.qe    = reg2hw.status_784.qe;
  assign rcache_line[3][16].status_reg.re    = reg2hw.status_784.re;


  assign rcache_line[3][17].tag_reg.tag      = reg2hw.tag_785.q;
  assign rcache_line[3][17].tag_reg.qe       = reg2hw.tag_785.qe;
  assign rcache_line[3][17].tag_reg.re       = reg2hw.tag_785.re;
  assign rcache_line[3][17].status_reg.status = reg2hw.status_785.q;//status_reg_t'(reg2hw.status_785.q);
  assign rcache_line[3][17].status_reg.qe    = reg2hw.status_785.qe;
  assign rcache_line[3][17].status_reg.re    = reg2hw.status_785.re;


  assign rcache_line[3][18].tag_reg.tag      = reg2hw.tag_786.q;
  assign rcache_line[3][18].tag_reg.qe       = reg2hw.tag_786.qe;
  assign rcache_line[3][18].tag_reg.re       = reg2hw.tag_786.re;
  assign rcache_line[3][18].status_reg.status = reg2hw.status_786.q;//status_reg_t'(reg2hw.status_786.q);
  assign rcache_line[3][18].status_reg.qe    = reg2hw.status_786.qe;
  assign rcache_line[3][18].status_reg.re    = reg2hw.status_786.re;


  assign rcache_line[3][19].tag_reg.tag      = reg2hw.tag_787.q;
  assign rcache_line[3][19].tag_reg.qe       = reg2hw.tag_787.qe;
  assign rcache_line[3][19].tag_reg.re       = reg2hw.tag_787.re;
  assign rcache_line[3][19].status_reg.status = reg2hw.status_787.q;//status_reg_t'(reg2hw.status_787.q);
  assign rcache_line[3][19].status_reg.qe    = reg2hw.status_787.qe;
  assign rcache_line[3][19].status_reg.re    = reg2hw.status_787.re;


  assign rcache_line[3][20].tag_reg.tag      = reg2hw.tag_788.q;
  assign rcache_line[3][20].tag_reg.qe       = reg2hw.tag_788.qe;
  assign rcache_line[3][20].tag_reg.re       = reg2hw.tag_788.re;
  assign rcache_line[3][20].status_reg.status = reg2hw.status_788.q;//status_reg_t'(reg2hw.status_788.q);
  assign rcache_line[3][20].status_reg.qe    = reg2hw.status_788.qe;
  assign rcache_line[3][20].status_reg.re    = reg2hw.status_788.re;


  assign rcache_line[3][21].tag_reg.tag      = reg2hw.tag_789.q;
  assign rcache_line[3][21].tag_reg.qe       = reg2hw.tag_789.qe;
  assign rcache_line[3][21].tag_reg.re       = reg2hw.tag_789.re;
  assign rcache_line[3][21].status_reg.status = reg2hw.status_789.q;//status_reg_t'(reg2hw.status_789.q);
  assign rcache_line[3][21].status_reg.qe    = reg2hw.status_789.qe;
  assign rcache_line[3][21].status_reg.re    = reg2hw.status_789.re;


  assign rcache_line[3][22].tag_reg.tag      = reg2hw.tag_790.q;
  assign rcache_line[3][22].tag_reg.qe       = reg2hw.tag_790.qe;
  assign rcache_line[3][22].tag_reg.re       = reg2hw.tag_790.re;
  assign rcache_line[3][22].status_reg.status = reg2hw.status_790.q;//status_reg_t'(reg2hw.status_790.q);
  assign rcache_line[3][22].status_reg.qe    = reg2hw.status_790.qe;
  assign rcache_line[3][22].status_reg.re    = reg2hw.status_790.re;


  assign rcache_line[3][23].tag_reg.tag      = reg2hw.tag_791.q;
  assign rcache_line[3][23].tag_reg.qe       = reg2hw.tag_791.qe;
  assign rcache_line[3][23].tag_reg.re       = reg2hw.tag_791.re;
  assign rcache_line[3][23].status_reg.status = reg2hw.status_791.q;//status_reg_t'(reg2hw.status_791.q);
  assign rcache_line[3][23].status_reg.qe    = reg2hw.status_791.qe;
  assign rcache_line[3][23].status_reg.re    = reg2hw.status_791.re;


  assign rcache_line[3][24].tag_reg.tag      = reg2hw.tag_792.q;
  assign rcache_line[3][24].tag_reg.qe       = reg2hw.tag_792.qe;
  assign rcache_line[3][24].tag_reg.re       = reg2hw.tag_792.re;
  assign rcache_line[3][24].status_reg.status = reg2hw.status_792.q;//status_reg_t'(reg2hw.status_792.q);
  assign rcache_line[3][24].status_reg.qe    = reg2hw.status_792.qe;
  assign rcache_line[3][24].status_reg.re    = reg2hw.status_792.re;


  assign rcache_line[3][25].tag_reg.tag      = reg2hw.tag_793.q;
  assign rcache_line[3][25].tag_reg.qe       = reg2hw.tag_793.qe;
  assign rcache_line[3][25].tag_reg.re       = reg2hw.tag_793.re;
  assign rcache_line[3][25].status_reg.status = reg2hw.status_793.q;//status_reg_t'(reg2hw.status_793.q);
  assign rcache_line[3][25].status_reg.qe    = reg2hw.status_793.qe;
  assign rcache_line[3][25].status_reg.re    = reg2hw.status_793.re;


  assign rcache_line[3][26].tag_reg.tag      = reg2hw.tag_794.q;
  assign rcache_line[3][26].tag_reg.qe       = reg2hw.tag_794.qe;
  assign rcache_line[3][26].tag_reg.re       = reg2hw.tag_794.re;
  assign rcache_line[3][26].status_reg.status = reg2hw.status_794.q;//status_reg_t'(reg2hw.status_794.q);
  assign rcache_line[3][26].status_reg.qe    = reg2hw.status_794.qe;
  assign rcache_line[3][26].status_reg.re    = reg2hw.status_794.re;


  assign rcache_line[3][27].tag_reg.tag      = reg2hw.tag_795.q;
  assign rcache_line[3][27].tag_reg.qe       = reg2hw.tag_795.qe;
  assign rcache_line[3][27].tag_reg.re       = reg2hw.tag_795.re;
  assign rcache_line[3][27].status_reg.status = reg2hw.status_795.q;//status_reg_t'(reg2hw.status_795.q);
  assign rcache_line[3][27].status_reg.qe    = reg2hw.status_795.qe;
  assign rcache_line[3][27].status_reg.re    = reg2hw.status_795.re;


  assign rcache_line[3][28].tag_reg.tag      = reg2hw.tag_796.q;
  assign rcache_line[3][28].tag_reg.qe       = reg2hw.tag_796.qe;
  assign rcache_line[3][28].tag_reg.re       = reg2hw.tag_796.re;
  assign rcache_line[3][28].status_reg.status = reg2hw.status_796.q;//status_reg_t'(reg2hw.status_796.q);
  assign rcache_line[3][28].status_reg.qe    = reg2hw.status_796.qe;
  assign rcache_line[3][28].status_reg.re    = reg2hw.status_796.re;


  assign rcache_line[3][29].tag_reg.tag      = reg2hw.tag_797.q;
  assign rcache_line[3][29].tag_reg.qe       = reg2hw.tag_797.qe;
  assign rcache_line[3][29].tag_reg.re       = reg2hw.tag_797.re;
  assign rcache_line[3][29].status_reg.status = reg2hw.status_797.q;//status_reg_t'(reg2hw.status_797.q);
  assign rcache_line[3][29].status_reg.qe    = reg2hw.status_797.qe;
  assign rcache_line[3][29].status_reg.re    = reg2hw.status_797.re;


  assign rcache_line[3][30].tag_reg.tag      = reg2hw.tag_798.q;
  assign rcache_line[3][30].tag_reg.qe       = reg2hw.tag_798.qe;
  assign rcache_line[3][30].tag_reg.re       = reg2hw.tag_798.re;
  assign rcache_line[3][30].status_reg.status = reg2hw.status_798.q;//status_reg_t'(reg2hw.status_798.q);
  assign rcache_line[3][30].status_reg.qe    = reg2hw.status_798.qe;
  assign rcache_line[3][30].status_reg.re    = reg2hw.status_798.re;


  assign rcache_line[3][31].tag_reg.tag      = reg2hw.tag_799.q;
  assign rcache_line[3][31].tag_reg.qe       = reg2hw.tag_799.qe;
  assign rcache_line[3][31].tag_reg.re       = reg2hw.tag_799.re;
  assign rcache_line[3][31].status_reg.status = reg2hw.status_799.q;//status_reg_t'(reg2hw.status_799.q);
  assign rcache_line[3][31].status_reg.qe    = reg2hw.status_799.qe;
  assign rcache_line[3][31].status_reg.re    = reg2hw.status_799.re;


  assign rcache_line[3][32].tag_reg.tag      = reg2hw.tag_800.q;
  assign rcache_line[3][32].tag_reg.qe       = reg2hw.tag_800.qe;
  assign rcache_line[3][32].tag_reg.re       = reg2hw.tag_800.re;
  assign rcache_line[3][32].status_reg.status = reg2hw.status_800.q;//status_reg_t'(reg2hw.status_800.q);
  assign rcache_line[3][32].status_reg.qe    = reg2hw.status_800.qe;
  assign rcache_line[3][32].status_reg.re    = reg2hw.status_800.re;


  assign rcache_line[3][33].tag_reg.tag      = reg2hw.tag_801.q;
  assign rcache_line[3][33].tag_reg.qe       = reg2hw.tag_801.qe;
  assign rcache_line[3][33].tag_reg.re       = reg2hw.tag_801.re;
  assign rcache_line[3][33].status_reg.status = reg2hw.status_801.q;//status_reg_t'(reg2hw.status_801.q);
  assign rcache_line[3][33].status_reg.qe    = reg2hw.status_801.qe;
  assign rcache_line[3][33].status_reg.re    = reg2hw.status_801.re;


  assign rcache_line[3][34].tag_reg.tag      = reg2hw.tag_802.q;
  assign rcache_line[3][34].tag_reg.qe       = reg2hw.tag_802.qe;
  assign rcache_line[3][34].tag_reg.re       = reg2hw.tag_802.re;
  assign rcache_line[3][34].status_reg.status = reg2hw.status_802.q;//status_reg_t'(reg2hw.status_802.q);
  assign rcache_line[3][34].status_reg.qe    = reg2hw.status_802.qe;
  assign rcache_line[3][34].status_reg.re    = reg2hw.status_802.re;


  assign rcache_line[3][35].tag_reg.tag      = reg2hw.tag_803.q;
  assign rcache_line[3][35].tag_reg.qe       = reg2hw.tag_803.qe;
  assign rcache_line[3][35].tag_reg.re       = reg2hw.tag_803.re;
  assign rcache_line[3][35].status_reg.status = reg2hw.status_803.q;//status_reg_t'(reg2hw.status_803.q);
  assign rcache_line[3][35].status_reg.qe    = reg2hw.status_803.qe;
  assign rcache_line[3][35].status_reg.re    = reg2hw.status_803.re;


  assign rcache_line[3][36].tag_reg.tag      = reg2hw.tag_804.q;
  assign rcache_line[3][36].tag_reg.qe       = reg2hw.tag_804.qe;
  assign rcache_line[3][36].tag_reg.re       = reg2hw.tag_804.re;
  assign rcache_line[3][36].status_reg.status = reg2hw.status_804.q;//status_reg_t'(reg2hw.status_804.q);
  assign rcache_line[3][36].status_reg.qe    = reg2hw.status_804.qe;
  assign rcache_line[3][36].status_reg.re    = reg2hw.status_804.re;


  assign rcache_line[3][37].tag_reg.tag      = reg2hw.tag_805.q;
  assign rcache_line[3][37].tag_reg.qe       = reg2hw.tag_805.qe;
  assign rcache_line[3][37].tag_reg.re       = reg2hw.tag_805.re;
  assign rcache_line[3][37].status_reg.status = reg2hw.status_805.q;//status_reg_t'(reg2hw.status_805.q);
  assign rcache_line[3][37].status_reg.qe    = reg2hw.status_805.qe;
  assign rcache_line[3][37].status_reg.re    = reg2hw.status_805.re;


  assign rcache_line[3][38].tag_reg.tag      = reg2hw.tag_806.q;
  assign rcache_line[3][38].tag_reg.qe       = reg2hw.tag_806.qe;
  assign rcache_line[3][38].tag_reg.re       = reg2hw.tag_806.re;
  assign rcache_line[3][38].status_reg.status = reg2hw.status_806.q;//status_reg_t'(reg2hw.status_806.q);
  assign rcache_line[3][38].status_reg.qe    = reg2hw.status_806.qe;
  assign rcache_line[3][38].status_reg.re    = reg2hw.status_806.re;


  assign rcache_line[3][39].tag_reg.tag      = reg2hw.tag_807.q;
  assign rcache_line[3][39].tag_reg.qe       = reg2hw.tag_807.qe;
  assign rcache_line[3][39].tag_reg.re       = reg2hw.tag_807.re;
  assign rcache_line[3][39].status_reg.status = reg2hw.status_807.q;//status_reg_t'(reg2hw.status_807.q);
  assign rcache_line[3][39].status_reg.qe    = reg2hw.status_807.qe;
  assign rcache_line[3][39].status_reg.re    = reg2hw.status_807.re;


  assign rcache_line[3][40].tag_reg.tag      = reg2hw.tag_808.q;
  assign rcache_line[3][40].tag_reg.qe       = reg2hw.tag_808.qe;
  assign rcache_line[3][40].tag_reg.re       = reg2hw.tag_808.re;
  assign rcache_line[3][40].status_reg.status = reg2hw.status_808.q;//status_reg_t'(reg2hw.status_808.q);
  assign rcache_line[3][40].status_reg.qe    = reg2hw.status_808.qe;
  assign rcache_line[3][40].status_reg.re    = reg2hw.status_808.re;


  assign rcache_line[3][41].tag_reg.tag      = reg2hw.tag_809.q;
  assign rcache_line[3][41].tag_reg.qe       = reg2hw.tag_809.qe;
  assign rcache_line[3][41].tag_reg.re       = reg2hw.tag_809.re;
  assign rcache_line[3][41].status_reg.status = reg2hw.status_809.q;//status_reg_t'(reg2hw.status_809.q);
  assign rcache_line[3][41].status_reg.qe    = reg2hw.status_809.qe;
  assign rcache_line[3][41].status_reg.re    = reg2hw.status_809.re;


  assign rcache_line[3][42].tag_reg.tag      = reg2hw.tag_810.q;
  assign rcache_line[3][42].tag_reg.qe       = reg2hw.tag_810.qe;
  assign rcache_line[3][42].tag_reg.re       = reg2hw.tag_810.re;
  assign rcache_line[3][42].status_reg.status = reg2hw.status_810.q;//status_reg_t'(reg2hw.status_810.q);
  assign rcache_line[3][42].status_reg.qe    = reg2hw.status_810.qe;
  assign rcache_line[3][42].status_reg.re    = reg2hw.status_810.re;


  assign rcache_line[3][43].tag_reg.tag      = reg2hw.tag_811.q;
  assign rcache_line[3][43].tag_reg.qe       = reg2hw.tag_811.qe;
  assign rcache_line[3][43].tag_reg.re       = reg2hw.tag_811.re;
  assign rcache_line[3][43].status_reg.status = reg2hw.status_811.q;//status_reg_t'(reg2hw.status_811.q);
  assign rcache_line[3][43].status_reg.qe    = reg2hw.status_811.qe;
  assign rcache_line[3][43].status_reg.re    = reg2hw.status_811.re;


  assign rcache_line[3][44].tag_reg.tag      = reg2hw.tag_812.q;
  assign rcache_line[3][44].tag_reg.qe       = reg2hw.tag_812.qe;
  assign rcache_line[3][44].tag_reg.re       = reg2hw.tag_812.re;
  assign rcache_line[3][44].status_reg.status = reg2hw.status_812.q;//status_reg_t'(reg2hw.status_812.q);
  assign rcache_line[3][44].status_reg.qe    = reg2hw.status_812.qe;
  assign rcache_line[3][44].status_reg.re    = reg2hw.status_812.re;


  assign rcache_line[3][45].tag_reg.tag      = reg2hw.tag_813.q;
  assign rcache_line[3][45].tag_reg.qe       = reg2hw.tag_813.qe;
  assign rcache_line[3][45].tag_reg.re       = reg2hw.tag_813.re;
  assign rcache_line[3][45].status_reg.status = reg2hw.status_813.q;//status_reg_t'(reg2hw.status_813.q);
  assign rcache_line[3][45].status_reg.qe    = reg2hw.status_813.qe;
  assign rcache_line[3][45].status_reg.re    = reg2hw.status_813.re;


  assign rcache_line[3][46].tag_reg.tag      = reg2hw.tag_814.q;
  assign rcache_line[3][46].tag_reg.qe       = reg2hw.tag_814.qe;
  assign rcache_line[3][46].tag_reg.re       = reg2hw.tag_814.re;
  assign rcache_line[3][46].status_reg.status = reg2hw.status_814.q;//status_reg_t'(reg2hw.status_814.q);
  assign rcache_line[3][46].status_reg.qe    = reg2hw.status_814.qe;
  assign rcache_line[3][46].status_reg.re    = reg2hw.status_814.re;


  assign rcache_line[3][47].tag_reg.tag      = reg2hw.tag_815.q;
  assign rcache_line[3][47].tag_reg.qe       = reg2hw.tag_815.qe;
  assign rcache_line[3][47].tag_reg.re       = reg2hw.tag_815.re;
  assign rcache_line[3][47].status_reg.status = reg2hw.status_815.q;//status_reg_t'(reg2hw.status_815.q);
  assign rcache_line[3][47].status_reg.qe    = reg2hw.status_815.qe;
  assign rcache_line[3][47].status_reg.re    = reg2hw.status_815.re;


  assign rcache_line[3][48].tag_reg.tag      = reg2hw.tag_816.q;
  assign rcache_line[3][48].tag_reg.qe       = reg2hw.tag_816.qe;
  assign rcache_line[3][48].tag_reg.re       = reg2hw.tag_816.re;
  assign rcache_line[3][48].status_reg.status = reg2hw.status_816.q;//status_reg_t'(reg2hw.status_816.q);
  assign rcache_line[3][48].status_reg.qe    = reg2hw.status_816.qe;
  assign rcache_line[3][48].status_reg.re    = reg2hw.status_816.re;


  assign rcache_line[3][49].tag_reg.tag      = reg2hw.tag_817.q;
  assign rcache_line[3][49].tag_reg.qe       = reg2hw.tag_817.qe;
  assign rcache_line[3][49].tag_reg.re       = reg2hw.tag_817.re;
  assign rcache_line[3][49].status_reg.status = reg2hw.status_817.q;//status_reg_t'(reg2hw.status_817.q);
  assign rcache_line[3][49].status_reg.qe    = reg2hw.status_817.qe;
  assign rcache_line[3][49].status_reg.re    = reg2hw.status_817.re;


  assign rcache_line[3][50].tag_reg.tag      = reg2hw.tag_818.q;
  assign rcache_line[3][50].tag_reg.qe       = reg2hw.tag_818.qe;
  assign rcache_line[3][50].tag_reg.re       = reg2hw.tag_818.re;
  assign rcache_line[3][50].status_reg.status = reg2hw.status_818.q;//status_reg_t'(reg2hw.status_818.q);
  assign rcache_line[3][50].status_reg.qe    = reg2hw.status_818.qe;
  assign rcache_line[3][50].status_reg.re    = reg2hw.status_818.re;


  assign rcache_line[3][51].tag_reg.tag      = reg2hw.tag_819.q;
  assign rcache_line[3][51].tag_reg.qe       = reg2hw.tag_819.qe;
  assign rcache_line[3][51].tag_reg.re       = reg2hw.tag_819.re;
  assign rcache_line[3][51].status_reg.status = reg2hw.status_819.q;//status_reg_t'(reg2hw.status_819.q);
  assign rcache_line[3][51].status_reg.qe    = reg2hw.status_819.qe;
  assign rcache_line[3][51].status_reg.re    = reg2hw.status_819.re;


  assign rcache_line[3][52].tag_reg.tag      = reg2hw.tag_820.q;
  assign rcache_line[3][52].tag_reg.qe       = reg2hw.tag_820.qe;
  assign rcache_line[3][52].tag_reg.re       = reg2hw.tag_820.re;
  assign rcache_line[3][52].status_reg.status = reg2hw.status_820.q;//status_reg_t'(reg2hw.status_820.q);
  assign rcache_line[3][52].status_reg.qe    = reg2hw.status_820.qe;
  assign rcache_line[3][52].status_reg.re    = reg2hw.status_820.re;


  assign rcache_line[3][53].tag_reg.tag      = reg2hw.tag_821.q;
  assign rcache_line[3][53].tag_reg.qe       = reg2hw.tag_821.qe;
  assign rcache_line[3][53].tag_reg.re       = reg2hw.tag_821.re;
  assign rcache_line[3][53].status_reg.status = reg2hw.status_821.q;//status_reg_t'(reg2hw.status_821.q);
  assign rcache_line[3][53].status_reg.qe    = reg2hw.status_821.qe;
  assign rcache_line[3][53].status_reg.re    = reg2hw.status_821.re;


  assign rcache_line[3][54].tag_reg.tag      = reg2hw.tag_822.q;
  assign rcache_line[3][54].tag_reg.qe       = reg2hw.tag_822.qe;
  assign rcache_line[3][54].tag_reg.re       = reg2hw.tag_822.re;
  assign rcache_line[3][54].status_reg.status = reg2hw.status_822.q;//status_reg_t'(reg2hw.status_822.q);
  assign rcache_line[3][54].status_reg.qe    = reg2hw.status_822.qe;
  assign rcache_line[3][54].status_reg.re    = reg2hw.status_822.re;


  assign rcache_line[3][55].tag_reg.tag      = reg2hw.tag_823.q;
  assign rcache_line[3][55].tag_reg.qe       = reg2hw.tag_823.qe;
  assign rcache_line[3][55].tag_reg.re       = reg2hw.tag_823.re;
  assign rcache_line[3][55].status_reg.status = reg2hw.status_823.q;//status_reg_t'(reg2hw.status_823.q);
  assign rcache_line[3][55].status_reg.qe    = reg2hw.status_823.qe;
  assign rcache_line[3][55].status_reg.re    = reg2hw.status_823.re;


  assign rcache_line[3][56].tag_reg.tag      = reg2hw.tag_824.q;
  assign rcache_line[3][56].tag_reg.qe       = reg2hw.tag_824.qe;
  assign rcache_line[3][56].tag_reg.re       = reg2hw.tag_824.re;
  assign rcache_line[3][56].status_reg.status = reg2hw.status_824.q;//status_reg_t'(reg2hw.status_824.q);
  assign rcache_line[3][56].status_reg.qe    = reg2hw.status_824.qe;
  assign rcache_line[3][56].status_reg.re    = reg2hw.status_824.re;


  assign rcache_line[3][57].tag_reg.tag      = reg2hw.tag_825.q;
  assign rcache_line[3][57].tag_reg.qe       = reg2hw.tag_825.qe;
  assign rcache_line[3][57].tag_reg.re       = reg2hw.tag_825.re;
  assign rcache_line[3][57].status_reg.status = reg2hw.status_825.q;//status_reg_t'(reg2hw.status_825.q);
  assign rcache_line[3][57].status_reg.qe    = reg2hw.status_825.qe;
  assign rcache_line[3][57].status_reg.re    = reg2hw.status_825.re;


  assign rcache_line[3][58].tag_reg.tag      = reg2hw.tag_826.q;
  assign rcache_line[3][58].tag_reg.qe       = reg2hw.tag_826.qe;
  assign rcache_line[3][58].tag_reg.re       = reg2hw.tag_826.re;
  assign rcache_line[3][58].status_reg.status = reg2hw.status_826.q;//status_reg_t'(reg2hw.status_826.q);
  assign rcache_line[3][58].status_reg.qe    = reg2hw.status_826.qe;
  assign rcache_line[3][58].status_reg.re    = reg2hw.status_826.re;


  assign rcache_line[3][59].tag_reg.tag      = reg2hw.tag_827.q;
  assign rcache_line[3][59].tag_reg.qe       = reg2hw.tag_827.qe;
  assign rcache_line[3][59].tag_reg.re       = reg2hw.tag_827.re;
  assign rcache_line[3][59].status_reg.status = reg2hw.status_827.q;//status_reg_t'(reg2hw.status_827.q);
  assign rcache_line[3][59].status_reg.qe    = reg2hw.status_827.qe;
  assign rcache_line[3][59].status_reg.re    = reg2hw.status_827.re;


  assign rcache_line[3][60].tag_reg.tag      = reg2hw.tag_828.q;
  assign rcache_line[3][60].tag_reg.qe       = reg2hw.tag_828.qe;
  assign rcache_line[3][60].tag_reg.re       = reg2hw.tag_828.re;
  assign rcache_line[3][60].status_reg.status = reg2hw.status_828.q;//status_reg_t'(reg2hw.status_828.q);
  assign rcache_line[3][60].status_reg.qe    = reg2hw.status_828.qe;
  assign rcache_line[3][60].status_reg.re    = reg2hw.status_828.re;


  assign rcache_line[3][61].tag_reg.tag      = reg2hw.tag_829.q;
  assign rcache_line[3][61].tag_reg.qe       = reg2hw.tag_829.qe;
  assign rcache_line[3][61].tag_reg.re       = reg2hw.tag_829.re;
  assign rcache_line[3][61].status_reg.status = reg2hw.status_829.q;//status_reg_t'(reg2hw.status_829.q);
  assign rcache_line[3][61].status_reg.qe    = reg2hw.status_829.qe;
  assign rcache_line[3][61].status_reg.re    = reg2hw.status_829.re;


  assign rcache_line[3][62].tag_reg.tag      = reg2hw.tag_830.q;
  assign rcache_line[3][62].tag_reg.qe       = reg2hw.tag_830.qe;
  assign rcache_line[3][62].tag_reg.re       = reg2hw.tag_830.re;
  assign rcache_line[3][62].status_reg.status = reg2hw.status_830.q;//status_reg_t'(reg2hw.status_830.q);
  assign rcache_line[3][62].status_reg.qe    = reg2hw.status_830.qe;
  assign rcache_line[3][62].status_reg.re    = reg2hw.status_830.re;


  assign rcache_line[3][63].tag_reg.tag      = reg2hw.tag_831.q;
  assign rcache_line[3][63].tag_reg.qe       = reg2hw.tag_831.qe;
  assign rcache_line[3][63].tag_reg.re       = reg2hw.tag_831.re;
  assign rcache_line[3][63].status_reg.status = reg2hw.status_831.q;//status_reg_t'(reg2hw.status_831.q);
  assign rcache_line[3][63].status_reg.qe    = reg2hw.status_831.qe;
  assign rcache_line[3][63].status_reg.re    = reg2hw.status_831.re;


  assign rcache_line[3][64].tag_reg.tag      = reg2hw.tag_832.q;
  assign rcache_line[3][64].tag_reg.qe       = reg2hw.tag_832.qe;
  assign rcache_line[3][64].tag_reg.re       = reg2hw.tag_832.re;
  assign rcache_line[3][64].status_reg.status = reg2hw.status_832.q;//status_reg_t'(reg2hw.status_832.q);
  assign rcache_line[3][64].status_reg.qe    = reg2hw.status_832.qe;
  assign rcache_line[3][64].status_reg.re    = reg2hw.status_832.re;


  assign rcache_line[3][65].tag_reg.tag      = reg2hw.tag_833.q;
  assign rcache_line[3][65].tag_reg.qe       = reg2hw.tag_833.qe;
  assign rcache_line[3][65].tag_reg.re       = reg2hw.tag_833.re;
  assign rcache_line[3][65].status_reg.status = reg2hw.status_833.q;//status_reg_t'(reg2hw.status_833.q);
  assign rcache_line[3][65].status_reg.qe    = reg2hw.status_833.qe;
  assign rcache_line[3][65].status_reg.re    = reg2hw.status_833.re;


  assign rcache_line[3][66].tag_reg.tag      = reg2hw.tag_834.q;
  assign rcache_line[3][66].tag_reg.qe       = reg2hw.tag_834.qe;
  assign rcache_line[3][66].tag_reg.re       = reg2hw.tag_834.re;
  assign rcache_line[3][66].status_reg.status = reg2hw.status_834.q;//status_reg_t'(reg2hw.status_834.q);
  assign rcache_line[3][66].status_reg.qe    = reg2hw.status_834.qe;
  assign rcache_line[3][66].status_reg.re    = reg2hw.status_834.re;


  assign rcache_line[3][67].tag_reg.tag      = reg2hw.tag_835.q;
  assign rcache_line[3][67].tag_reg.qe       = reg2hw.tag_835.qe;
  assign rcache_line[3][67].tag_reg.re       = reg2hw.tag_835.re;
  assign rcache_line[3][67].status_reg.status = reg2hw.status_835.q;//status_reg_t'(reg2hw.status_835.q);
  assign rcache_line[3][67].status_reg.qe    = reg2hw.status_835.qe;
  assign rcache_line[3][67].status_reg.re    = reg2hw.status_835.re;


  assign rcache_line[3][68].tag_reg.tag      = reg2hw.tag_836.q;
  assign rcache_line[3][68].tag_reg.qe       = reg2hw.tag_836.qe;
  assign rcache_line[3][68].tag_reg.re       = reg2hw.tag_836.re;
  assign rcache_line[3][68].status_reg.status = reg2hw.status_836.q;//status_reg_t'(reg2hw.status_836.q);
  assign rcache_line[3][68].status_reg.qe    = reg2hw.status_836.qe;
  assign rcache_line[3][68].status_reg.re    = reg2hw.status_836.re;


  assign rcache_line[3][69].tag_reg.tag      = reg2hw.tag_837.q;
  assign rcache_line[3][69].tag_reg.qe       = reg2hw.tag_837.qe;
  assign rcache_line[3][69].tag_reg.re       = reg2hw.tag_837.re;
  assign rcache_line[3][69].status_reg.status = reg2hw.status_837.q;//status_reg_t'(reg2hw.status_837.q);
  assign rcache_line[3][69].status_reg.qe    = reg2hw.status_837.qe;
  assign rcache_line[3][69].status_reg.re    = reg2hw.status_837.re;


  assign rcache_line[3][70].tag_reg.tag      = reg2hw.tag_838.q;
  assign rcache_line[3][70].tag_reg.qe       = reg2hw.tag_838.qe;
  assign rcache_line[3][70].tag_reg.re       = reg2hw.tag_838.re;
  assign rcache_line[3][70].status_reg.status = reg2hw.status_838.q;//status_reg_t'(reg2hw.status_838.q);
  assign rcache_line[3][70].status_reg.qe    = reg2hw.status_838.qe;
  assign rcache_line[3][70].status_reg.re    = reg2hw.status_838.re;


  assign rcache_line[3][71].tag_reg.tag      = reg2hw.tag_839.q;
  assign rcache_line[3][71].tag_reg.qe       = reg2hw.tag_839.qe;
  assign rcache_line[3][71].tag_reg.re       = reg2hw.tag_839.re;
  assign rcache_line[3][71].status_reg.status = reg2hw.status_839.q;//status_reg_t'(reg2hw.status_839.q);
  assign rcache_line[3][71].status_reg.qe    = reg2hw.status_839.qe;
  assign rcache_line[3][71].status_reg.re    = reg2hw.status_839.re;


  assign rcache_line[3][72].tag_reg.tag      = reg2hw.tag_840.q;
  assign rcache_line[3][72].tag_reg.qe       = reg2hw.tag_840.qe;
  assign rcache_line[3][72].tag_reg.re       = reg2hw.tag_840.re;
  assign rcache_line[3][72].status_reg.status = reg2hw.status_840.q;//status_reg_t'(reg2hw.status_840.q);
  assign rcache_line[3][72].status_reg.qe    = reg2hw.status_840.qe;
  assign rcache_line[3][72].status_reg.re    = reg2hw.status_840.re;


  assign rcache_line[3][73].tag_reg.tag      = reg2hw.tag_841.q;
  assign rcache_line[3][73].tag_reg.qe       = reg2hw.tag_841.qe;
  assign rcache_line[3][73].tag_reg.re       = reg2hw.tag_841.re;
  assign rcache_line[3][73].status_reg.status = reg2hw.status_841.q;//status_reg_t'(reg2hw.status_841.q);
  assign rcache_line[3][73].status_reg.qe    = reg2hw.status_841.qe;
  assign rcache_line[3][73].status_reg.re    = reg2hw.status_841.re;


  assign rcache_line[3][74].tag_reg.tag      = reg2hw.tag_842.q;
  assign rcache_line[3][74].tag_reg.qe       = reg2hw.tag_842.qe;
  assign rcache_line[3][74].tag_reg.re       = reg2hw.tag_842.re;
  assign rcache_line[3][74].status_reg.status = reg2hw.status_842.q;//status_reg_t'(reg2hw.status_842.q);
  assign rcache_line[3][74].status_reg.qe    = reg2hw.status_842.qe;
  assign rcache_line[3][74].status_reg.re    = reg2hw.status_842.re;


  assign rcache_line[3][75].tag_reg.tag      = reg2hw.tag_843.q;
  assign rcache_line[3][75].tag_reg.qe       = reg2hw.tag_843.qe;
  assign rcache_line[3][75].tag_reg.re       = reg2hw.tag_843.re;
  assign rcache_line[3][75].status_reg.status = reg2hw.status_843.q;//status_reg_t'(reg2hw.status_843.q);
  assign rcache_line[3][75].status_reg.qe    = reg2hw.status_843.qe;
  assign rcache_line[3][75].status_reg.re    = reg2hw.status_843.re;


  assign rcache_line[3][76].tag_reg.tag      = reg2hw.tag_844.q;
  assign rcache_line[3][76].tag_reg.qe       = reg2hw.tag_844.qe;
  assign rcache_line[3][76].tag_reg.re       = reg2hw.tag_844.re;
  assign rcache_line[3][76].status_reg.status = reg2hw.status_844.q;//status_reg_t'(reg2hw.status_844.q);
  assign rcache_line[3][76].status_reg.qe    = reg2hw.status_844.qe;
  assign rcache_line[3][76].status_reg.re    = reg2hw.status_844.re;


  assign rcache_line[3][77].tag_reg.tag      = reg2hw.tag_845.q;
  assign rcache_line[3][77].tag_reg.qe       = reg2hw.tag_845.qe;
  assign rcache_line[3][77].tag_reg.re       = reg2hw.tag_845.re;
  assign rcache_line[3][77].status_reg.status = reg2hw.status_845.q;//status_reg_t'(reg2hw.status_845.q);
  assign rcache_line[3][77].status_reg.qe    = reg2hw.status_845.qe;
  assign rcache_line[3][77].status_reg.re    = reg2hw.status_845.re;


  assign rcache_line[3][78].tag_reg.tag      = reg2hw.tag_846.q;
  assign rcache_line[3][78].tag_reg.qe       = reg2hw.tag_846.qe;
  assign rcache_line[3][78].tag_reg.re       = reg2hw.tag_846.re;
  assign rcache_line[3][78].status_reg.status = reg2hw.status_846.q;//status_reg_t'(reg2hw.status_846.q);
  assign rcache_line[3][78].status_reg.qe    = reg2hw.status_846.qe;
  assign rcache_line[3][78].status_reg.re    = reg2hw.status_846.re;


  assign rcache_line[3][79].tag_reg.tag      = reg2hw.tag_847.q;
  assign rcache_line[3][79].tag_reg.qe       = reg2hw.tag_847.qe;
  assign rcache_line[3][79].tag_reg.re       = reg2hw.tag_847.re;
  assign rcache_line[3][79].status_reg.status = reg2hw.status_847.q;//status_reg_t'(reg2hw.status_847.q);
  assign rcache_line[3][79].status_reg.qe    = reg2hw.status_847.qe;
  assign rcache_line[3][79].status_reg.re    = reg2hw.status_847.re;


  assign rcache_line[3][80].tag_reg.tag      = reg2hw.tag_848.q;
  assign rcache_line[3][80].tag_reg.qe       = reg2hw.tag_848.qe;
  assign rcache_line[3][80].tag_reg.re       = reg2hw.tag_848.re;
  assign rcache_line[3][80].status_reg.status = reg2hw.status_848.q;//status_reg_t'(reg2hw.status_848.q);
  assign rcache_line[3][80].status_reg.qe    = reg2hw.status_848.qe;
  assign rcache_line[3][80].status_reg.re    = reg2hw.status_848.re;


  assign rcache_line[3][81].tag_reg.tag      = reg2hw.tag_849.q;
  assign rcache_line[3][81].tag_reg.qe       = reg2hw.tag_849.qe;
  assign rcache_line[3][81].tag_reg.re       = reg2hw.tag_849.re;
  assign rcache_line[3][81].status_reg.status = reg2hw.status_849.q;//status_reg_t'(reg2hw.status_849.q);
  assign rcache_line[3][81].status_reg.qe    = reg2hw.status_849.qe;
  assign rcache_line[3][81].status_reg.re    = reg2hw.status_849.re;


  assign rcache_line[3][82].tag_reg.tag      = reg2hw.tag_850.q;
  assign rcache_line[3][82].tag_reg.qe       = reg2hw.tag_850.qe;
  assign rcache_line[3][82].tag_reg.re       = reg2hw.tag_850.re;
  assign rcache_line[3][82].status_reg.status = reg2hw.status_850.q;//status_reg_t'(reg2hw.status_850.q);
  assign rcache_line[3][82].status_reg.qe    = reg2hw.status_850.qe;
  assign rcache_line[3][82].status_reg.re    = reg2hw.status_850.re;


  assign rcache_line[3][83].tag_reg.tag      = reg2hw.tag_851.q;
  assign rcache_line[3][83].tag_reg.qe       = reg2hw.tag_851.qe;
  assign rcache_line[3][83].tag_reg.re       = reg2hw.tag_851.re;
  assign rcache_line[3][83].status_reg.status = reg2hw.status_851.q;//status_reg_t'(reg2hw.status_851.q);
  assign rcache_line[3][83].status_reg.qe    = reg2hw.status_851.qe;
  assign rcache_line[3][83].status_reg.re    = reg2hw.status_851.re;


  assign rcache_line[3][84].tag_reg.tag      = reg2hw.tag_852.q;
  assign rcache_line[3][84].tag_reg.qe       = reg2hw.tag_852.qe;
  assign rcache_line[3][84].tag_reg.re       = reg2hw.tag_852.re;
  assign rcache_line[3][84].status_reg.status = reg2hw.status_852.q;//status_reg_t'(reg2hw.status_852.q);
  assign rcache_line[3][84].status_reg.qe    = reg2hw.status_852.qe;
  assign rcache_line[3][84].status_reg.re    = reg2hw.status_852.re;


  assign rcache_line[3][85].tag_reg.tag      = reg2hw.tag_853.q;
  assign rcache_line[3][85].tag_reg.qe       = reg2hw.tag_853.qe;
  assign rcache_line[3][85].tag_reg.re       = reg2hw.tag_853.re;
  assign rcache_line[3][85].status_reg.status = reg2hw.status_853.q;//status_reg_t'(reg2hw.status_853.q);
  assign rcache_line[3][85].status_reg.qe    = reg2hw.status_853.qe;
  assign rcache_line[3][85].status_reg.re    = reg2hw.status_853.re;


  assign rcache_line[3][86].tag_reg.tag      = reg2hw.tag_854.q;
  assign rcache_line[3][86].tag_reg.qe       = reg2hw.tag_854.qe;
  assign rcache_line[3][86].tag_reg.re       = reg2hw.tag_854.re;
  assign rcache_line[3][86].status_reg.status = reg2hw.status_854.q;//status_reg_t'(reg2hw.status_854.q);
  assign rcache_line[3][86].status_reg.qe    = reg2hw.status_854.qe;
  assign rcache_line[3][86].status_reg.re    = reg2hw.status_854.re;


  assign rcache_line[3][87].tag_reg.tag      = reg2hw.tag_855.q;
  assign rcache_line[3][87].tag_reg.qe       = reg2hw.tag_855.qe;
  assign rcache_line[3][87].tag_reg.re       = reg2hw.tag_855.re;
  assign rcache_line[3][87].status_reg.status = reg2hw.status_855.q;//status_reg_t'(reg2hw.status_855.q);
  assign rcache_line[3][87].status_reg.qe    = reg2hw.status_855.qe;
  assign rcache_line[3][87].status_reg.re    = reg2hw.status_855.re;


  assign rcache_line[3][88].tag_reg.tag      = reg2hw.tag_856.q;
  assign rcache_line[3][88].tag_reg.qe       = reg2hw.tag_856.qe;
  assign rcache_line[3][88].tag_reg.re       = reg2hw.tag_856.re;
  assign rcache_line[3][88].status_reg.status = reg2hw.status_856.q;//status_reg_t'(reg2hw.status_856.q);
  assign rcache_line[3][88].status_reg.qe    = reg2hw.status_856.qe;
  assign rcache_line[3][88].status_reg.re    = reg2hw.status_856.re;


  assign rcache_line[3][89].tag_reg.tag      = reg2hw.tag_857.q;
  assign rcache_line[3][89].tag_reg.qe       = reg2hw.tag_857.qe;
  assign rcache_line[3][89].tag_reg.re       = reg2hw.tag_857.re;
  assign rcache_line[3][89].status_reg.status = reg2hw.status_857.q;//status_reg_t'(reg2hw.status_857.q);
  assign rcache_line[3][89].status_reg.qe    = reg2hw.status_857.qe;
  assign rcache_line[3][89].status_reg.re    = reg2hw.status_857.re;


  assign rcache_line[3][90].tag_reg.tag      = reg2hw.tag_858.q;
  assign rcache_line[3][90].tag_reg.qe       = reg2hw.tag_858.qe;
  assign rcache_line[3][90].tag_reg.re       = reg2hw.tag_858.re;
  assign rcache_line[3][90].status_reg.status = reg2hw.status_858.q;//status_reg_t'(reg2hw.status_858.q);
  assign rcache_line[3][90].status_reg.qe    = reg2hw.status_858.qe;
  assign rcache_line[3][90].status_reg.re    = reg2hw.status_858.re;


  assign rcache_line[3][91].tag_reg.tag      = reg2hw.tag_859.q;
  assign rcache_line[3][91].tag_reg.qe       = reg2hw.tag_859.qe;
  assign rcache_line[3][91].tag_reg.re       = reg2hw.tag_859.re;
  assign rcache_line[3][91].status_reg.status = reg2hw.status_859.q;//status_reg_t'(reg2hw.status_859.q);
  assign rcache_line[3][91].status_reg.qe    = reg2hw.status_859.qe;
  assign rcache_line[3][91].status_reg.re    = reg2hw.status_859.re;


  assign rcache_line[3][92].tag_reg.tag      = reg2hw.tag_860.q;
  assign rcache_line[3][92].tag_reg.qe       = reg2hw.tag_860.qe;
  assign rcache_line[3][92].tag_reg.re       = reg2hw.tag_860.re;
  assign rcache_line[3][92].status_reg.status = reg2hw.status_860.q;//status_reg_t'(reg2hw.status_860.q);
  assign rcache_line[3][92].status_reg.qe    = reg2hw.status_860.qe;
  assign rcache_line[3][92].status_reg.re    = reg2hw.status_860.re;


  assign rcache_line[3][93].tag_reg.tag      = reg2hw.tag_861.q;
  assign rcache_line[3][93].tag_reg.qe       = reg2hw.tag_861.qe;
  assign rcache_line[3][93].tag_reg.re       = reg2hw.tag_861.re;
  assign rcache_line[3][93].status_reg.status = reg2hw.status_861.q;//status_reg_t'(reg2hw.status_861.q);
  assign rcache_line[3][93].status_reg.qe    = reg2hw.status_861.qe;
  assign rcache_line[3][93].status_reg.re    = reg2hw.status_861.re;


  assign rcache_line[3][94].tag_reg.tag      = reg2hw.tag_862.q;
  assign rcache_line[3][94].tag_reg.qe       = reg2hw.tag_862.qe;
  assign rcache_line[3][94].tag_reg.re       = reg2hw.tag_862.re;
  assign rcache_line[3][94].status_reg.status = reg2hw.status_862.q;//status_reg_t'(reg2hw.status_862.q);
  assign rcache_line[3][94].status_reg.qe    = reg2hw.status_862.qe;
  assign rcache_line[3][94].status_reg.re    = reg2hw.status_862.re;


  assign rcache_line[3][95].tag_reg.tag      = reg2hw.tag_863.q;
  assign rcache_line[3][95].tag_reg.qe       = reg2hw.tag_863.qe;
  assign rcache_line[3][95].tag_reg.re       = reg2hw.tag_863.re;
  assign rcache_line[3][95].status_reg.status = reg2hw.status_863.q;//status_reg_t'(reg2hw.status_863.q);
  assign rcache_line[3][95].status_reg.qe    = reg2hw.status_863.qe;
  assign rcache_line[3][95].status_reg.re    = reg2hw.status_863.re;


  assign rcache_line[3][96].tag_reg.tag      = reg2hw.tag_864.q;
  assign rcache_line[3][96].tag_reg.qe       = reg2hw.tag_864.qe;
  assign rcache_line[3][96].tag_reg.re       = reg2hw.tag_864.re;
  assign rcache_line[3][96].status_reg.status = reg2hw.status_864.q;//status_reg_t'(reg2hw.status_864.q);
  assign rcache_line[3][96].status_reg.qe    = reg2hw.status_864.qe;
  assign rcache_line[3][96].status_reg.re    = reg2hw.status_864.re;


  assign rcache_line[3][97].tag_reg.tag      = reg2hw.tag_865.q;
  assign rcache_line[3][97].tag_reg.qe       = reg2hw.tag_865.qe;
  assign rcache_line[3][97].tag_reg.re       = reg2hw.tag_865.re;
  assign rcache_line[3][97].status_reg.status = reg2hw.status_865.q;//status_reg_t'(reg2hw.status_865.q);
  assign rcache_line[3][97].status_reg.qe    = reg2hw.status_865.qe;
  assign rcache_line[3][97].status_reg.re    = reg2hw.status_865.re;


  assign rcache_line[3][98].tag_reg.tag      = reg2hw.tag_866.q;
  assign rcache_line[3][98].tag_reg.qe       = reg2hw.tag_866.qe;
  assign rcache_line[3][98].tag_reg.re       = reg2hw.tag_866.re;
  assign rcache_line[3][98].status_reg.status = reg2hw.status_866.q;//status_reg_t'(reg2hw.status_866.q);
  assign rcache_line[3][98].status_reg.qe    = reg2hw.status_866.qe;
  assign rcache_line[3][98].status_reg.re    = reg2hw.status_866.re;


  assign rcache_line[3][99].tag_reg.tag      = reg2hw.tag_867.q;
  assign rcache_line[3][99].tag_reg.qe       = reg2hw.tag_867.qe;
  assign rcache_line[3][99].tag_reg.re       = reg2hw.tag_867.re;
  assign rcache_line[3][99].status_reg.status = reg2hw.status_867.q;//status_reg_t'(reg2hw.status_867.q);
  assign rcache_line[3][99].status_reg.qe    = reg2hw.status_867.qe;
  assign rcache_line[3][99].status_reg.re    = reg2hw.status_867.re;


  assign rcache_line[3][100].tag_reg.tag      = reg2hw.tag_868.q;
  assign rcache_line[3][100].tag_reg.qe       = reg2hw.tag_868.qe;
  assign rcache_line[3][100].tag_reg.re       = reg2hw.tag_868.re;
  assign rcache_line[3][100].status_reg.status = reg2hw.status_868.q;//status_reg_t'(reg2hw.status_868.q);
  assign rcache_line[3][100].status_reg.qe    = reg2hw.status_868.qe;
  assign rcache_line[3][100].status_reg.re    = reg2hw.status_868.re;


  assign rcache_line[3][101].tag_reg.tag      = reg2hw.tag_869.q;
  assign rcache_line[3][101].tag_reg.qe       = reg2hw.tag_869.qe;
  assign rcache_line[3][101].tag_reg.re       = reg2hw.tag_869.re;
  assign rcache_line[3][101].status_reg.status = reg2hw.status_869.q;//status_reg_t'(reg2hw.status_869.q);
  assign rcache_line[3][101].status_reg.qe    = reg2hw.status_869.qe;
  assign rcache_line[3][101].status_reg.re    = reg2hw.status_869.re;


  assign rcache_line[3][102].tag_reg.tag      = reg2hw.tag_870.q;
  assign rcache_line[3][102].tag_reg.qe       = reg2hw.tag_870.qe;
  assign rcache_line[3][102].tag_reg.re       = reg2hw.tag_870.re;
  assign rcache_line[3][102].status_reg.status = reg2hw.status_870.q;//status_reg_t'(reg2hw.status_870.q);
  assign rcache_line[3][102].status_reg.qe    = reg2hw.status_870.qe;
  assign rcache_line[3][102].status_reg.re    = reg2hw.status_870.re;


  assign rcache_line[3][103].tag_reg.tag      = reg2hw.tag_871.q;
  assign rcache_line[3][103].tag_reg.qe       = reg2hw.tag_871.qe;
  assign rcache_line[3][103].tag_reg.re       = reg2hw.tag_871.re;
  assign rcache_line[3][103].status_reg.status = reg2hw.status_871.q;//status_reg_t'(reg2hw.status_871.q);
  assign rcache_line[3][103].status_reg.qe    = reg2hw.status_871.qe;
  assign rcache_line[3][103].status_reg.re    = reg2hw.status_871.re;


  assign rcache_line[3][104].tag_reg.tag      = reg2hw.tag_872.q;
  assign rcache_line[3][104].tag_reg.qe       = reg2hw.tag_872.qe;
  assign rcache_line[3][104].tag_reg.re       = reg2hw.tag_872.re;
  assign rcache_line[3][104].status_reg.status = reg2hw.status_872.q;//status_reg_t'(reg2hw.status_872.q);
  assign rcache_line[3][104].status_reg.qe    = reg2hw.status_872.qe;
  assign rcache_line[3][104].status_reg.re    = reg2hw.status_872.re;


  assign rcache_line[3][105].tag_reg.tag      = reg2hw.tag_873.q;
  assign rcache_line[3][105].tag_reg.qe       = reg2hw.tag_873.qe;
  assign rcache_line[3][105].tag_reg.re       = reg2hw.tag_873.re;
  assign rcache_line[3][105].status_reg.status = reg2hw.status_873.q;//status_reg_t'(reg2hw.status_873.q);
  assign rcache_line[3][105].status_reg.qe    = reg2hw.status_873.qe;
  assign rcache_line[3][105].status_reg.re    = reg2hw.status_873.re;


  assign rcache_line[3][106].tag_reg.tag      = reg2hw.tag_874.q;
  assign rcache_line[3][106].tag_reg.qe       = reg2hw.tag_874.qe;
  assign rcache_line[3][106].tag_reg.re       = reg2hw.tag_874.re;
  assign rcache_line[3][106].status_reg.status = reg2hw.status_874.q;//status_reg_t'(reg2hw.status_874.q);
  assign rcache_line[3][106].status_reg.qe    = reg2hw.status_874.qe;
  assign rcache_line[3][106].status_reg.re    = reg2hw.status_874.re;


  assign rcache_line[3][107].tag_reg.tag      = reg2hw.tag_875.q;
  assign rcache_line[3][107].tag_reg.qe       = reg2hw.tag_875.qe;
  assign rcache_line[3][107].tag_reg.re       = reg2hw.tag_875.re;
  assign rcache_line[3][107].status_reg.status = reg2hw.status_875.q;//status_reg_t'(reg2hw.status_875.q);
  assign rcache_line[3][107].status_reg.qe    = reg2hw.status_875.qe;
  assign rcache_line[3][107].status_reg.re    = reg2hw.status_875.re;


  assign rcache_line[3][108].tag_reg.tag      = reg2hw.tag_876.q;
  assign rcache_line[3][108].tag_reg.qe       = reg2hw.tag_876.qe;
  assign rcache_line[3][108].tag_reg.re       = reg2hw.tag_876.re;
  assign rcache_line[3][108].status_reg.status = reg2hw.status_876.q;//status_reg_t'(reg2hw.status_876.q);
  assign rcache_line[3][108].status_reg.qe    = reg2hw.status_876.qe;
  assign rcache_line[3][108].status_reg.re    = reg2hw.status_876.re;


  assign rcache_line[3][109].tag_reg.tag      = reg2hw.tag_877.q;
  assign rcache_line[3][109].tag_reg.qe       = reg2hw.tag_877.qe;
  assign rcache_line[3][109].tag_reg.re       = reg2hw.tag_877.re;
  assign rcache_line[3][109].status_reg.status = reg2hw.status_877.q;//status_reg_t'(reg2hw.status_877.q);
  assign rcache_line[3][109].status_reg.qe    = reg2hw.status_877.qe;
  assign rcache_line[3][109].status_reg.re    = reg2hw.status_877.re;


  assign rcache_line[3][110].tag_reg.tag      = reg2hw.tag_878.q;
  assign rcache_line[3][110].tag_reg.qe       = reg2hw.tag_878.qe;
  assign rcache_line[3][110].tag_reg.re       = reg2hw.tag_878.re;
  assign rcache_line[3][110].status_reg.status = reg2hw.status_878.q;//status_reg_t'(reg2hw.status_878.q);
  assign rcache_line[3][110].status_reg.qe    = reg2hw.status_878.qe;
  assign rcache_line[3][110].status_reg.re    = reg2hw.status_878.re;


  assign rcache_line[3][111].tag_reg.tag      = reg2hw.tag_879.q;
  assign rcache_line[3][111].tag_reg.qe       = reg2hw.tag_879.qe;
  assign rcache_line[3][111].tag_reg.re       = reg2hw.tag_879.re;
  assign rcache_line[3][111].status_reg.status = reg2hw.status_879.q;//status_reg_t'(reg2hw.status_879.q);
  assign rcache_line[3][111].status_reg.qe    = reg2hw.status_879.qe;
  assign rcache_line[3][111].status_reg.re    = reg2hw.status_879.re;


  assign rcache_line[3][112].tag_reg.tag      = reg2hw.tag_880.q;
  assign rcache_line[3][112].tag_reg.qe       = reg2hw.tag_880.qe;
  assign rcache_line[3][112].tag_reg.re       = reg2hw.tag_880.re;
  assign rcache_line[3][112].status_reg.status = reg2hw.status_880.q;//status_reg_t'(reg2hw.status_880.q);
  assign rcache_line[3][112].status_reg.qe    = reg2hw.status_880.qe;
  assign rcache_line[3][112].status_reg.re    = reg2hw.status_880.re;


  assign rcache_line[3][113].tag_reg.tag      = reg2hw.tag_881.q;
  assign rcache_line[3][113].tag_reg.qe       = reg2hw.tag_881.qe;
  assign rcache_line[3][113].tag_reg.re       = reg2hw.tag_881.re;
  assign rcache_line[3][113].status_reg.status = reg2hw.status_881.q;//status_reg_t'(reg2hw.status_881.q);
  assign rcache_line[3][113].status_reg.qe    = reg2hw.status_881.qe;
  assign rcache_line[3][113].status_reg.re    = reg2hw.status_881.re;


  assign rcache_line[3][114].tag_reg.tag      = reg2hw.tag_882.q;
  assign rcache_line[3][114].tag_reg.qe       = reg2hw.tag_882.qe;
  assign rcache_line[3][114].tag_reg.re       = reg2hw.tag_882.re;
  assign rcache_line[3][114].status_reg.status = reg2hw.status_882.q;//status_reg_t'(reg2hw.status_882.q);
  assign rcache_line[3][114].status_reg.qe    = reg2hw.status_882.qe;
  assign rcache_line[3][114].status_reg.re    = reg2hw.status_882.re;


  assign rcache_line[3][115].tag_reg.tag      = reg2hw.tag_883.q;
  assign rcache_line[3][115].tag_reg.qe       = reg2hw.tag_883.qe;
  assign rcache_line[3][115].tag_reg.re       = reg2hw.tag_883.re;
  assign rcache_line[3][115].status_reg.status = reg2hw.status_883.q;//status_reg_t'(reg2hw.status_883.q);
  assign rcache_line[3][115].status_reg.qe    = reg2hw.status_883.qe;
  assign rcache_line[3][115].status_reg.re    = reg2hw.status_883.re;


  assign rcache_line[3][116].tag_reg.tag      = reg2hw.tag_884.q;
  assign rcache_line[3][116].tag_reg.qe       = reg2hw.tag_884.qe;
  assign rcache_line[3][116].tag_reg.re       = reg2hw.tag_884.re;
  assign rcache_line[3][116].status_reg.status = reg2hw.status_884.q;//status_reg_t'(reg2hw.status_884.q);
  assign rcache_line[3][116].status_reg.qe    = reg2hw.status_884.qe;
  assign rcache_line[3][116].status_reg.re    = reg2hw.status_884.re;


  assign rcache_line[3][117].tag_reg.tag      = reg2hw.tag_885.q;
  assign rcache_line[3][117].tag_reg.qe       = reg2hw.tag_885.qe;
  assign rcache_line[3][117].tag_reg.re       = reg2hw.tag_885.re;
  assign rcache_line[3][117].status_reg.status = reg2hw.status_885.q;//status_reg_t'(reg2hw.status_885.q);
  assign rcache_line[3][117].status_reg.qe    = reg2hw.status_885.qe;
  assign rcache_line[3][117].status_reg.re    = reg2hw.status_885.re;


  assign rcache_line[3][118].tag_reg.tag      = reg2hw.tag_886.q;
  assign rcache_line[3][118].tag_reg.qe       = reg2hw.tag_886.qe;
  assign rcache_line[3][118].tag_reg.re       = reg2hw.tag_886.re;
  assign rcache_line[3][118].status_reg.status = reg2hw.status_886.q;//status_reg_t'(reg2hw.status_886.q);
  assign rcache_line[3][118].status_reg.qe    = reg2hw.status_886.qe;
  assign rcache_line[3][118].status_reg.re    = reg2hw.status_886.re;


  assign rcache_line[3][119].tag_reg.tag      = reg2hw.tag_887.q;
  assign rcache_line[3][119].tag_reg.qe       = reg2hw.tag_887.qe;
  assign rcache_line[3][119].tag_reg.re       = reg2hw.tag_887.re;
  assign rcache_line[3][119].status_reg.status = reg2hw.status_887.q;//status_reg_t'(reg2hw.status_887.q);
  assign rcache_line[3][119].status_reg.qe    = reg2hw.status_887.qe;
  assign rcache_line[3][119].status_reg.re    = reg2hw.status_887.re;


  assign rcache_line[3][120].tag_reg.tag      = reg2hw.tag_888.q;
  assign rcache_line[3][120].tag_reg.qe       = reg2hw.tag_888.qe;
  assign rcache_line[3][120].tag_reg.re       = reg2hw.tag_888.re;
  assign rcache_line[3][120].status_reg.status = reg2hw.status_888.q;//status_reg_t'(reg2hw.status_888.q);
  assign rcache_line[3][120].status_reg.qe    = reg2hw.status_888.qe;
  assign rcache_line[3][120].status_reg.re    = reg2hw.status_888.re;


  assign rcache_line[3][121].tag_reg.tag      = reg2hw.tag_889.q;
  assign rcache_line[3][121].tag_reg.qe       = reg2hw.tag_889.qe;
  assign rcache_line[3][121].tag_reg.re       = reg2hw.tag_889.re;
  assign rcache_line[3][121].status_reg.status = reg2hw.status_889.q;//status_reg_t'(reg2hw.status_889.q);
  assign rcache_line[3][121].status_reg.qe    = reg2hw.status_889.qe;
  assign rcache_line[3][121].status_reg.re    = reg2hw.status_889.re;


  assign rcache_line[3][122].tag_reg.tag      = reg2hw.tag_890.q;
  assign rcache_line[3][122].tag_reg.qe       = reg2hw.tag_890.qe;
  assign rcache_line[3][122].tag_reg.re       = reg2hw.tag_890.re;
  assign rcache_line[3][122].status_reg.status = reg2hw.status_890.q;//status_reg_t'(reg2hw.status_890.q);
  assign rcache_line[3][122].status_reg.qe    = reg2hw.status_890.qe;
  assign rcache_line[3][122].status_reg.re    = reg2hw.status_890.re;


  assign rcache_line[3][123].tag_reg.tag      = reg2hw.tag_891.q;
  assign rcache_line[3][123].tag_reg.qe       = reg2hw.tag_891.qe;
  assign rcache_line[3][123].tag_reg.re       = reg2hw.tag_891.re;
  assign rcache_line[3][123].status_reg.status = reg2hw.status_891.q;//status_reg_t'(reg2hw.status_891.q);
  assign rcache_line[3][123].status_reg.qe    = reg2hw.status_891.qe;
  assign rcache_line[3][123].status_reg.re    = reg2hw.status_891.re;


  assign rcache_line[3][124].tag_reg.tag      = reg2hw.tag_892.q;
  assign rcache_line[3][124].tag_reg.qe       = reg2hw.tag_892.qe;
  assign rcache_line[3][124].tag_reg.re       = reg2hw.tag_892.re;
  assign rcache_line[3][124].status_reg.status = reg2hw.status_892.q;//status_reg_t'(reg2hw.status_892.q);
  assign rcache_line[3][124].status_reg.qe    = reg2hw.status_892.qe;
  assign rcache_line[3][124].status_reg.re    = reg2hw.status_892.re;


  assign rcache_line[3][125].tag_reg.tag      = reg2hw.tag_893.q;
  assign rcache_line[3][125].tag_reg.qe       = reg2hw.tag_893.qe;
  assign rcache_line[3][125].tag_reg.re       = reg2hw.tag_893.re;
  assign rcache_line[3][125].status_reg.status = reg2hw.status_893.q;//status_reg_t'(reg2hw.status_893.q);
  assign rcache_line[3][125].status_reg.qe    = reg2hw.status_893.qe;
  assign rcache_line[3][125].status_reg.re    = reg2hw.status_893.re;


  assign rcache_line[3][126].tag_reg.tag      = reg2hw.tag_894.q;
  assign rcache_line[3][126].tag_reg.qe       = reg2hw.tag_894.qe;
  assign rcache_line[3][126].tag_reg.re       = reg2hw.tag_894.re;
  assign rcache_line[3][126].status_reg.status = reg2hw.status_894.q;//status_reg_t'(reg2hw.status_894.q);
  assign rcache_line[3][126].status_reg.qe    = reg2hw.status_894.qe;
  assign rcache_line[3][126].status_reg.re    = reg2hw.status_894.re;


  assign rcache_line[3][127].tag_reg.tag      = reg2hw.tag_895.q;
  assign rcache_line[3][127].tag_reg.qe       = reg2hw.tag_895.qe;
  assign rcache_line[3][127].tag_reg.re       = reg2hw.tag_895.re;
  assign rcache_line[3][127].status_reg.status = reg2hw.status_895.q;//status_reg_t'(reg2hw.status_895.q);
  assign rcache_line[3][127].status_reg.qe    = reg2hw.status_895.qe;
  assign rcache_line[3][127].status_reg.re    = reg2hw.status_895.re;


  assign rcache_line[3][128].tag_reg.tag      = reg2hw.tag_896.q;
  assign rcache_line[3][128].tag_reg.qe       = reg2hw.tag_896.qe;
  assign rcache_line[3][128].tag_reg.re       = reg2hw.tag_896.re;
  assign rcache_line[3][128].status_reg.status = reg2hw.status_896.q;//status_reg_t'(reg2hw.status_896.q);
  assign rcache_line[3][128].status_reg.qe    = reg2hw.status_896.qe;
  assign rcache_line[3][128].status_reg.re    = reg2hw.status_896.re;


  assign rcache_line[3][129].tag_reg.tag      = reg2hw.tag_897.q;
  assign rcache_line[3][129].tag_reg.qe       = reg2hw.tag_897.qe;
  assign rcache_line[3][129].tag_reg.re       = reg2hw.tag_897.re;
  assign rcache_line[3][129].status_reg.status = reg2hw.status_897.q;//status_reg_t'(reg2hw.status_897.q);
  assign rcache_line[3][129].status_reg.qe    = reg2hw.status_897.qe;
  assign rcache_line[3][129].status_reg.re    = reg2hw.status_897.re;


  assign rcache_line[3][130].tag_reg.tag      = reg2hw.tag_898.q;
  assign rcache_line[3][130].tag_reg.qe       = reg2hw.tag_898.qe;
  assign rcache_line[3][130].tag_reg.re       = reg2hw.tag_898.re;
  assign rcache_line[3][130].status_reg.status = reg2hw.status_898.q;//status_reg_t'(reg2hw.status_898.q);
  assign rcache_line[3][130].status_reg.qe    = reg2hw.status_898.qe;
  assign rcache_line[3][130].status_reg.re    = reg2hw.status_898.re;


  assign rcache_line[3][131].tag_reg.tag      = reg2hw.tag_899.q;
  assign rcache_line[3][131].tag_reg.qe       = reg2hw.tag_899.qe;
  assign rcache_line[3][131].tag_reg.re       = reg2hw.tag_899.re;
  assign rcache_line[3][131].status_reg.status = reg2hw.status_899.q;//status_reg_t'(reg2hw.status_899.q);
  assign rcache_line[3][131].status_reg.qe    = reg2hw.status_899.qe;
  assign rcache_line[3][131].status_reg.re    = reg2hw.status_899.re;


  assign rcache_line[3][132].tag_reg.tag      = reg2hw.tag_900.q;
  assign rcache_line[3][132].tag_reg.qe       = reg2hw.tag_900.qe;
  assign rcache_line[3][132].tag_reg.re       = reg2hw.tag_900.re;
  assign rcache_line[3][132].status_reg.status = reg2hw.status_900.q;//status_reg_t'(reg2hw.status_900.q);
  assign rcache_line[3][132].status_reg.qe    = reg2hw.status_900.qe;
  assign rcache_line[3][132].status_reg.re    = reg2hw.status_900.re;


  assign rcache_line[3][133].tag_reg.tag      = reg2hw.tag_901.q;
  assign rcache_line[3][133].tag_reg.qe       = reg2hw.tag_901.qe;
  assign rcache_line[3][133].tag_reg.re       = reg2hw.tag_901.re;
  assign rcache_line[3][133].status_reg.status = reg2hw.status_901.q;//status_reg_t'(reg2hw.status_901.q);
  assign rcache_line[3][133].status_reg.qe    = reg2hw.status_901.qe;
  assign rcache_line[3][133].status_reg.re    = reg2hw.status_901.re;


  assign rcache_line[3][134].tag_reg.tag      = reg2hw.tag_902.q;
  assign rcache_line[3][134].tag_reg.qe       = reg2hw.tag_902.qe;
  assign rcache_line[3][134].tag_reg.re       = reg2hw.tag_902.re;
  assign rcache_line[3][134].status_reg.status = reg2hw.status_902.q;//status_reg_t'(reg2hw.status_902.q);
  assign rcache_line[3][134].status_reg.qe    = reg2hw.status_902.qe;
  assign rcache_line[3][134].status_reg.re    = reg2hw.status_902.re;


  assign rcache_line[3][135].tag_reg.tag      = reg2hw.tag_903.q;
  assign rcache_line[3][135].tag_reg.qe       = reg2hw.tag_903.qe;
  assign rcache_line[3][135].tag_reg.re       = reg2hw.tag_903.re;
  assign rcache_line[3][135].status_reg.status = reg2hw.status_903.q;//status_reg_t'(reg2hw.status_903.q);
  assign rcache_line[3][135].status_reg.qe    = reg2hw.status_903.qe;
  assign rcache_line[3][135].status_reg.re    = reg2hw.status_903.re;


  assign rcache_line[3][136].tag_reg.tag      = reg2hw.tag_904.q;
  assign rcache_line[3][136].tag_reg.qe       = reg2hw.tag_904.qe;
  assign rcache_line[3][136].tag_reg.re       = reg2hw.tag_904.re;
  assign rcache_line[3][136].status_reg.status = reg2hw.status_904.q;//status_reg_t'(reg2hw.status_904.q);
  assign rcache_line[3][136].status_reg.qe    = reg2hw.status_904.qe;
  assign rcache_line[3][136].status_reg.re    = reg2hw.status_904.re;


  assign rcache_line[3][137].tag_reg.tag      = reg2hw.tag_905.q;
  assign rcache_line[3][137].tag_reg.qe       = reg2hw.tag_905.qe;
  assign rcache_line[3][137].tag_reg.re       = reg2hw.tag_905.re;
  assign rcache_line[3][137].status_reg.status = reg2hw.status_905.q;//status_reg_t'(reg2hw.status_905.q);
  assign rcache_line[3][137].status_reg.qe    = reg2hw.status_905.qe;
  assign rcache_line[3][137].status_reg.re    = reg2hw.status_905.re;


  assign rcache_line[3][138].tag_reg.tag      = reg2hw.tag_906.q;
  assign rcache_line[3][138].tag_reg.qe       = reg2hw.tag_906.qe;
  assign rcache_line[3][138].tag_reg.re       = reg2hw.tag_906.re;
  assign rcache_line[3][138].status_reg.status = reg2hw.status_906.q;//status_reg_t'(reg2hw.status_906.q);
  assign rcache_line[3][138].status_reg.qe    = reg2hw.status_906.qe;
  assign rcache_line[3][138].status_reg.re    = reg2hw.status_906.re;


  assign rcache_line[3][139].tag_reg.tag      = reg2hw.tag_907.q;
  assign rcache_line[3][139].tag_reg.qe       = reg2hw.tag_907.qe;
  assign rcache_line[3][139].tag_reg.re       = reg2hw.tag_907.re;
  assign rcache_line[3][139].status_reg.status = reg2hw.status_907.q;//status_reg_t'(reg2hw.status_907.q);
  assign rcache_line[3][139].status_reg.qe    = reg2hw.status_907.qe;
  assign rcache_line[3][139].status_reg.re    = reg2hw.status_907.re;


  assign rcache_line[3][140].tag_reg.tag      = reg2hw.tag_908.q;
  assign rcache_line[3][140].tag_reg.qe       = reg2hw.tag_908.qe;
  assign rcache_line[3][140].tag_reg.re       = reg2hw.tag_908.re;
  assign rcache_line[3][140].status_reg.status = reg2hw.status_908.q;//status_reg_t'(reg2hw.status_908.q);
  assign rcache_line[3][140].status_reg.qe    = reg2hw.status_908.qe;
  assign rcache_line[3][140].status_reg.re    = reg2hw.status_908.re;


  assign rcache_line[3][141].tag_reg.tag      = reg2hw.tag_909.q;
  assign rcache_line[3][141].tag_reg.qe       = reg2hw.tag_909.qe;
  assign rcache_line[3][141].tag_reg.re       = reg2hw.tag_909.re;
  assign rcache_line[3][141].status_reg.status = reg2hw.status_909.q;//status_reg_t'(reg2hw.status_909.q);
  assign rcache_line[3][141].status_reg.qe    = reg2hw.status_909.qe;
  assign rcache_line[3][141].status_reg.re    = reg2hw.status_909.re;


  assign rcache_line[3][142].tag_reg.tag      = reg2hw.tag_910.q;
  assign rcache_line[3][142].tag_reg.qe       = reg2hw.tag_910.qe;
  assign rcache_line[3][142].tag_reg.re       = reg2hw.tag_910.re;
  assign rcache_line[3][142].status_reg.status = reg2hw.status_910.q;//status_reg_t'(reg2hw.status_910.q);
  assign rcache_line[3][142].status_reg.qe    = reg2hw.status_910.qe;
  assign rcache_line[3][142].status_reg.re    = reg2hw.status_910.re;


  assign rcache_line[3][143].tag_reg.tag      = reg2hw.tag_911.q;
  assign rcache_line[3][143].tag_reg.qe       = reg2hw.tag_911.qe;
  assign rcache_line[3][143].tag_reg.re       = reg2hw.tag_911.re;
  assign rcache_line[3][143].status_reg.status = reg2hw.status_911.q;//status_reg_t'(reg2hw.status_911.q);
  assign rcache_line[3][143].status_reg.qe    = reg2hw.status_911.qe;
  assign rcache_line[3][143].status_reg.re    = reg2hw.status_911.re;


  assign rcache_line[3][144].tag_reg.tag      = reg2hw.tag_912.q;
  assign rcache_line[3][144].tag_reg.qe       = reg2hw.tag_912.qe;
  assign rcache_line[3][144].tag_reg.re       = reg2hw.tag_912.re;
  assign rcache_line[3][144].status_reg.status = reg2hw.status_912.q;//status_reg_t'(reg2hw.status_912.q);
  assign rcache_line[3][144].status_reg.qe    = reg2hw.status_912.qe;
  assign rcache_line[3][144].status_reg.re    = reg2hw.status_912.re;


  assign rcache_line[3][145].tag_reg.tag      = reg2hw.tag_913.q;
  assign rcache_line[3][145].tag_reg.qe       = reg2hw.tag_913.qe;
  assign rcache_line[3][145].tag_reg.re       = reg2hw.tag_913.re;
  assign rcache_line[3][145].status_reg.status = reg2hw.status_913.q;//status_reg_t'(reg2hw.status_913.q);
  assign rcache_line[3][145].status_reg.qe    = reg2hw.status_913.qe;
  assign rcache_line[3][145].status_reg.re    = reg2hw.status_913.re;


  assign rcache_line[3][146].tag_reg.tag      = reg2hw.tag_914.q;
  assign rcache_line[3][146].tag_reg.qe       = reg2hw.tag_914.qe;
  assign rcache_line[3][146].tag_reg.re       = reg2hw.tag_914.re;
  assign rcache_line[3][146].status_reg.status = reg2hw.status_914.q;//status_reg_t'(reg2hw.status_914.q);
  assign rcache_line[3][146].status_reg.qe    = reg2hw.status_914.qe;
  assign rcache_line[3][146].status_reg.re    = reg2hw.status_914.re;


  assign rcache_line[3][147].tag_reg.tag      = reg2hw.tag_915.q;
  assign rcache_line[3][147].tag_reg.qe       = reg2hw.tag_915.qe;
  assign rcache_line[3][147].tag_reg.re       = reg2hw.tag_915.re;
  assign rcache_line[3][147].status_reg.status = reg2hw.status_915.q;//status_reg_t'(reg2hw.status_915.q);
  assign rcache_line[3][147].status_reg.qe    = reg2hw.status_915.qe;
  assign rcache_line[3][147].status_reg.re    = reg2hw.status_915.re;


  assign rcache_line[3][148].tag_reg.tag      = reg2hw.tag_916.q;
  assign rcache_line[3][148].tag_reg.qe       = reg2hw.tag_916.qe;
  assign rcache_line[3][148].tag_reg.re       = reg2hw.tag_916.re;
  assign rcache_line[3][148].status_reg.status = reg2hw.status_916.q;//status_reg_t'(reg2hw.status_916.q);
  assign rcache_line[3][148].status_reg.qe    = reg2hw.status_916.qe;
  assign rcache_line[3][148].status_reg.re    = reg2hw.status_916.re;


  assign rcache_line[3][149].tag_reg.tag      = reg2hw.tag_917.q;
  assign rcache_line[3][149].tag_reg.qe       = reg2hw.tag_917.qe;
  assign rcache_line[3][149].tag_reg.re       = reg2hw.tag_917.re;
  assign rcache_line[3][149].status_reg.status = reg2hw.status_917.q;//status_reg_t'(reg2hw.status_917.q);
  assign rcache_line[3][149].status_reg.qe    = reg2hw.status_917.qe;
  assign rcache_line[3][149].status_reg.re    = reg2hw.status_917.re;


  assign rcache_line[3][150].tag_reg.tag      = reg2hw.tag_918.q;
  assign rcache_line[3][150].tag_reg.qe       = reg2hw.tag_918.qe;
  assign rcache_line[3][150].tag_reg.re       = reg2hw.tag_918.re;
  assign rcache_line[3][150].status_reg.status = reg2hw.status_918.q;//status_reg_t'(reg2hw.status_918.q);
  assign rcache_line[3][150].status_reg.qe    = reg2hw.status_918.qe;
  assign rcache_line[3][150].status_reg.re    = reg2hw.status_918.re;


  assign rcache_line[3][151].tag_reg.tag      = reg2hw.tag_919.q;
  assign rcache_line[3][151].tag_reg.qe       = reg2hw.tag_919.qe;
  assign rcache_line[3][151].tag_reg.re       = reg2hw.tag_919.re;
  assign rcache_line[3][151].status_reg.status = reg2hw.status_919.q;//status_reg_t'(reg2hw.status_919.q);
  assign rcache_line[3][151].status_reg.qe    = reg2hw.status_919.qe;
  assign rcache_line[3][151].status_reg.re    = reg2hw.status_919.re;


  assign rcache_line[3][152].tag_reg.tag      = reg2hw.tag_920.q;
  assign rcache_line[3][152].tag_reg.qe       = reg2hw.tag_920.qe;
  assign rcache_line[3][152].tag_reg.re       = reg2hw.tag_920.re;
  assign rcache_line[3][152].status_reg.status = reg2hw.status_920.q;//status_reg_t'(reg2hw.status_920.q);
  assign rcache_line[3][152].status_reg.qe    = reg2hw.status_920.qe;
  assign rcache_line[3][152].status_reg.re    = reg2hw.status_920.re;


  assign rcache_line[3][153].tag_reg.tag      = reg2hw.tag_921.q;
  assign rcache_line[3][153].tag_reg.qe       = reg2hw.tag_921.qe;
  assign rcache_line[3][153].tag_reg.re       = reg2hw.tag_921.re;
  assign rcache_line[3][153].status_reg.status = reg2hw.status_921.q;//status_reg_t'(reg2hw.status_921.q);
  assign rcache_line[3][153].status_reg.qe    = reg2hw.status_921.qe;
  assign rcache_line[3][153].status_reg.re    = reg2hw.status_921.re;


  assign rcache_line[3][154].tag_reg.tag      = reg2hw.tag_922.q;
  assign rcache_line[3][154].tag_reg.qe       = reg2hw.tag_922.qe;
  assign rcache_line[3][154].tag_reg.re       = reg2hw.tag_922.re;
  assign rcache_line[3][154].status_reg.status = reg2hw.status_922.q;//status_reg_t'(reg2hw.status_922.q);
  assign rcache_line[3][154].status_reg.qe    = reg2hw.status_922.qe;
  assign rcache_line[3][154].status_reg.re    = reg2hw.status_922.re;


  assign rcache_line[3][155].tag_reg.tag      = reg2hw.tag_923.q;
  assign rcache_line[3][155].tag_reg.qe       = reg2hw.tag_923.qe;
  assign rcache_line[3][155].tag_reg.re       = reg2hw.tag_923.re;
  assign rcache_line[3][155].status_reg.status = reg2hw.status_923.q;//status_reg_t'(reg2hw.status_923.q);
  assign rcache_line[3][155].status_reg.qe    = reg2hw.status_923.qe;
  assign rcache_line[3][155].status_reg.re    = reg2hw.status_923.re;


  assign rcache_line[3][156].tag_reg.tag      = reg2hw.tag_924.q;
  assign rcache_line[3][156].tag_reg.qe       = reg2hw.tag_924.qe;
  assign rcache_line[3][156].tag_reg.re       = reg2hw.tag_924.re;
  assign rcache_line[3][156].status_reg.status = reg2hw.status_924.q;//status_reg_t'(reg2hw.status_924.q);
  assign rcache_line[3][156].status_reg.qe    = reg2hw.status_924.qe;
  assign rcache_line[3][156].status_reg.re    = reg2hw.status_924.re;


  assign rcache_line[3][157].tag_reg.tag      = reg2hw.tag_925.q;
  assign rcache_line[3][157].tag_reg.qe       = reg2hw.tag_925.qe;
  assign rcache_line[3][157].tag_reg.re       = reg2hw.tag_925.re;
  assign rcache_line[3][157].status_reg.status = reg2hw.status_925.q;//status_reg_t'(reg2hw.status_925.q);
  assign rcache_line[3][157].status_reg.qe    = reg2hw.status_925.qe;
  assign rcache_line[3][157].status_reg.re    = reg2hw.status_925.re;


  assign rcache_line[3][158].tag_reg.tag      = reg2hw.tag_926.q;
  assign rcache_line[3][158].tag_reg.qe       = reg2hw.tag_926.qe;
  assign rcache_line[3][158].tag_reg.re       = reg2hw.tag_926.re;
  assign rcache_line[3][158].status_reg.status = reg2hw.status_926.q;//status_reg_t'(reg2hw.status_926.q);
  assign rcache_line[3][158].status_reg.qe    = reg2hw.status_926.qe;
  assign rcache_line[3][158].status_reg.re    = reg2hw.status_926.re;


  assign rcache_line[3][159].tag_reg.tag      = reg2hw.tag_927.q;
  assign rcache_line[3][159].tag_reg.qe       = reg2hw.tag_927.qe;
  assign rcache_line[3][159].tag_reg.re       = reg2hw.tag_927.re;
  assign rcache_line[3][159].status_reg.status = reg2hw.status_927.q;//status_reg_t'(reg2hw.status_927.q);
  assign rcache_line[3][159].status_reg.qe    = reg2hw.status_927.qe;
  assign rcache_line[3][159].status_reg.re    = reg2hw.status_927.re;


  assign rcache_line[3][160].tag_reg.tag      = reg2hw.tag_928.q;
  assign rcache_line[3][160].tag_reg.qe       = reg2hw.tag_928.qe;
  assign rcache_line[3][160].tag_reg.re       = reg2hw.tag_928.re;
  assign rcache_line[3][160].status_reg.status = reg2hw.status_928.q;//status_reg_t'(reg2hw.status_928.q);
  assign rcache_line[3][160].status_reg.qe    = reg2hw.status_928.qe;
  assign rcache_line[3][160].status_reg.re    = reg2hw.status_928.re;


  assign rcache_line[3][161].tag_reg.tag      = reg2hw.tag_929.q;
  assign rcache_line[3][161].tag_reg.qe       = reg2hw.tag_929.qe;
  assign rcache_line[3][161].tag_reg.re       = reg2hw.tag_929.re;
  assign rcache_line[3][161].status_reg.status = reg2hw.status_929.q;//status_reg_t'(reg2hw.status_929.q);
  assign rcache_line[3][161].status_reg.qe    = reg2hw.status_929.qe;
  assign rcache_line[3][161].status_reg.re    = reg2hw.status_929.re;


  assign rcache_line[3][162].tag_reg.tag      = reg2hw.tag_930.q;
  assign rcache_line[3][162].tag_reg.qe       = reg2hw.tag_930.qe;
  assign rcache_line[3][162].tag_reg.re       = reg2hw.tag_930.re;
  assign rcache_line[3][162].status_reg.status = reg2hw.status_930.q;//status_reg_t'(reg2hw.status_930.q);
  assign rcache_line[3][162].status_reg.qe    = reg2hw.status_930.qe;
  assign rcache_line[3][162].status_reg.re    = reg2hw.status_930.re;


  assign rcache_line[3][163].tag_reg.tag      = reg2hw.tag_931.q;
  assign rcache_line[3][163].tag_reg.qe       = reg2hw.tag_931.qe;
  assign rcache_line[3][163].tag_reg.re       = reg2hw.tag_931.re;
  assign rcache_line[3][163].status_reg.status = reg2hw.status_931.q;//status_reg_t'(reg2hw.status_931.q);
  assign rcache_line[3][163].status_reg.qe    = reg2hw.status_931.qe;
  assign rcache_line[3][163].status_reg.re    = reg2hw.status_931.re;


  assign rcache_line[3][164].tag_reg.tag      = reg2hw.tag_932.q;
  assign rcache_line[3][164].tag_reg.qe       = reg2hw.tag_932.qe;
  assign rcache_line[3][164].tag_reg.re       = reg2hw.tag_932.re;
  assign rcache_line[3][164].status_reg.status = reg2hw.status_932.q;//status_reg_t'(reg2hw.status_932.q);
  assign rcache_line[3][164].status_reg.qe    = reg2hw.status_932.qe;
  assign rcache_line[3][164].status_reg.re    = reg2hw.status_932.re;


  assign rcache_line[3][165].tag_reg.tag      = reg2hw.tag_933.q;
  assign rcache_line[3][165].tag_reg.qe       = reg2hw.tag_933.qe;
  assign rcache_line[3][165].tag_reg.re       = reg2hw.tag_933.re;
  assign rcache_line[3][165].status_reg.status = reg2hw.status_933.q;//status_reg_t'(reg2hw.status_933.q);
  assign rcache_line[3][165].status_reg.qe    = reg2hw.status_933.qe;
  assign rcache_line[3][165].status_reg.re    = reg2hw.status_933.re;


  assign rcache_line[3][166].tag_reg.tag      = reg2hw.tag_934.q;
  assign rcache_line[3][166].tag_reg.qe       = reg2hw.tag_934.qe;
  assign rcache_line[3][166].tag_reg.re       = reg2hw.tag_934.re;
  assign rcache_line[3][166].status_reg.status = reg2hw.status_934.q;//status_reg_t'(reg2hw.status_934.q);
  assign rcache_line[3][166].status_reg.qe    = reg2hw.status_934.qe;
  assign rcache_line[3][166].status_reg.re    = reg2hw.status_934.re;


  assign rcache_line[3][167].tag_reg.tag      = reg2hw.tag_935.q;
  assign rcache_line[3][167].tag_reg.qe       = reg2hw.tag_935.qe;
  assign rcache_line[3][167].tag_reg.re       = reg2hw.tag_935.re;
  assign rcache_line[3][167].status_reg.status = reg2hw.status_935.q;//status_reg_t'(reg2hw.status_935.q);
  assign rcache_line[3][167].status_reg.qe    = reg2hw.status_935.qe;
  assign rcache_line[3][167].status_reg.re    = reg2hw.status_935.re;


  assign rcache_line[3][168].tag_reg.tag      = reg2hw.tag_936.q;
  assign rcache_line[3][168].tag_reg.qe       = reg2hw.tag_936.qe;
  assign rcache_line[3][168].tag_reg.re       = reg2hw.tag_936.re;
  assign rcache_line[3][168].status_reg.status = reg2hw.status_936.q;//status_reg_t'(reg2hw.status_936.q);
  assign rcache_line[3][168].status_reg.qe    = reg2hw.status_936.qe;
  assign rcache_line[3][168].status_reg.re    = reg2hw.status_936.re;


  assign rcache_line[3][169].tag_reg.tag      = reg2hw.tag_937.q;
  assign rcache_line[3][169].tag_reg.qe       = reg2hw.tag_937.qe;
  assign rcache_line[3][169].tag_reg.re       = reg2hw.tag_937.re;
  assign rcache_line[3][169].status_reg.status = reg2hw.status_937.q;//status_reg_t'(reg2hw.status_937.q);
  assign rcache_line[3][169].status_reg.qe    = reg2hw.status_937.qe;
  assign rcache_line[3][169].status_reg.re    = reg2hw.status_937.re;


  assign rcache_line[3][170].tag_reg.tag      = reg2hw.tag_938.q;
  assign rcache_line[3][170].tag_reg.qe       = reg2hw.tag_938.qe;
  assign rcache_line[3][170].tag_reg.re       = reg2hw.tag_938.re;
  assign rcache_line[3][170].status_reg.status = reg2hw.status_938.q;//status_reg_t'(reg2hw.status_938.q);
  assign rcache_line[3][170].status_reg.qe    = reg2hw.status_938.qe;
  assign rcache_line[3][170].status_reg.re    = reg2hw.status_938.re;


  assign rcache_line[3][171].tag_reg.tag      = reg2hw.tag_939.q;
  assign rcache_line[3][171].tag_reg.qe       = reg2hw.tag_939.qe;
  assign rcache_line[3][171].tag_reg.re       = reg2hw.tag_939.re;
  assign rcache_line[3][171].status_reg.status = reg2hw.status_939.q;//status_reg_t'(reg2hw.status_939.q);
  assign rcache_line[3][171].status_reg.qe    = reg2hw.status_939.qe;
  assign rcache_line[3][171].status_reg.re    = reg2hw.status_939.re;


  assign rcache_line[3][172].tag_reg.tag      = reg2hw.tag_940.q;
  assign rcache_line[3][172].tag_reg.qe       = reg2hw.tag_940.qe;
  assign rcache_line[3][172].tag_reg.re       = reg2hw.tag_940.re;
  assign rcache_line[3][172].status_reg.status = reg2hw.status_940.q;//status_reg_t'(reg2hw.status_940.q);
  assign rcache_line[3][172].status_reg.qe    = reg2hw.status_940.qe;
  assign rcache_line[3][172].status_reg.re    = reg2hw.status_940.re;


  assign rcache_line[3][173].tag_reg.tag      = reg2hw.tag_941.q;
  assign rcache_line[3][173].tag_reg.qe       = reg2hw.tag_941.qe;
  assign rcache_line[3][173].tag_reg.re       = reg2hw.tag_941.re;
  assign rcache_line[3][173].status_reg.status = reg2hw.status_941.q;//status_reg_t'(reg2hw.status_941.q);
  assign rcache_line[3][173].status_reg.qe    = reg2hw.status_941.qe;
  assign rcache_line[3][173].status_reg.re    = reg2hw.status_941.re;


  assign rcache_line[3][174].tag_reg.tag      = reg2hw.tag_942.q;
  assign rcache_line[3][174].tag_reg.qe       = reg2hw.tag_942.qe;
  assign rcache_line[3][174].tag_reg.re       = reg2hw.tag_942.re;
  assign rcache_line[3][174].status_reg.status = reg2hw.status_942.q;//status_reg_t'(reg2hw.status_942.q);
  assign rcache_line[3][174].status_reg.qe    = reg2hw.status_942.qe;
  assign rcache_line[3][174].status_reg.re    = reg2hw.status_942.re;


  assign rcache_line[3][175].tag_reg.tag      = reg2hw.tag_943.q;
  assign rcache_line[3][175].tag_reg.qe       = reg2hw.tag_943.qe;
  assign rcache_line[3][175].tag_reg.re       = reg2hw.tag_943.re;
  assign rcache_line[3][175].status_reg.status = reg2hw.status_943.q;//status_reg_t'(reg2hw.status_943.q);
  assign rcache_line[3][175].status_reg.qe    = reg2hw.status_943.qe;
  assign rcache_line[3][175].status_reg.re    = reg2hw.status_943.re;


  assign rcache_line[3][176].tag_reg.tag      = reg2hw.tag_944.q;
  assign rcache_line[3][176].tag_reg.qe       = reg2hw.tag_944.qe;
  assign rcache_line[3][176].tag_reg.re       = reg2hw.tag_944.re;
  assign rcache_line[3][176].status_reg.status = reg2hw.status_944.q;//status_reg_t'(reg2hw.status_944.q);
  assign rcache_line[3][176].status_reg.qe    = reg2hw.status_944.qe;
  assign rcache_line[3][176].status_reg.re    = reg2hw.status_944.re;


  assign rcache_line[3][177].tag_reg.tag      = reg2hw.tag_945.q;
  assign rcache_line[3][177].tag_reg.qe       = reg2hw.tag_945.qe;
  assign rcache_line[3][177].tag_reg.re       = reg2hw.tag_945.re;
  assign rcache_line[3][177].status_reg.status = reg2hw.status_945.q;//status_reg_t'(reg2hw.status_945.q);
  assign rcache_line[3][177].status_reg.qe    = reg2hw.status_945.qe;
  assign rcache_line[3][177].status_reg.re    = reg2hw.status_945.re;


  assign rcache_line[3][178].tag_reg.tag      = reg2hw.tag_946.q;
  assign rcache_line[3][178].tag_reg.qe       = reg2hw.tag_946.qe;
  assign rcache_line[3][178].tag_reg.re       = reg2hw.tag_946.re;
  assign rcache_line[3][178].status_reg.status = reg2hw.status_946.q;//status_reg_t'(reg2hw.status_946.q);
  assign rcache_line[3][178].status_reg.qe    = reg2hw.status_946.qe;
  assign rcache_line[3][178].status_reg.re    = reg2hw.status_946.re;


  assign rcache_line[3][179].tag_reg.tag      = reg2hw.tag_947.q;
  assign rcache_line[3][179].tag_reg.qe       = reg2hw.tag_947.qe;
  assign rcache_line[3][179].tag_reg.re       = reg2hw.tag_947.re;
  assign rcache_line[3][179].status_reg.status = reg2hw.status_947.q;//status_reg_t'(reg2hw.status_947.q);
  assign rcache_line[3][179].status_reg.qe    = reg2hw.status_947.qe;
  assign rcache_line[3][179].status_reg.re    = reg2hw.status_947.re;


  assign rcache_line[3][180].tag_reg.tag      = reg2hw.tag_948.q;
  assign rcache_line[3][180].tag_reg.qe       = reg2hw.tag_948.qe;
  assign rcache_line[3][180].tag_reg.re       = reg2hw.tag_948.re;
  assign rcache_line[3][180].status_reg.status = reg2hw.status_948.q;//status_reg_t'(reg2hw.status_948.q);
  assign rcache_line[3][180].status_reg.qe    = reg2hw.status_948.qe;
  assign rcache_line[3][180].status_reg.re    = reg2hw.status_948.re;


  assign rcache_line[3][181].tag_reg.tag      = reg2hw.tag_949.q;
  assign rcache_line[3][181].tag_reg.qe       = reg2hw.tag_949.qe;
  assign rcache_line[3][181].tag_reg.re       = reg2hw.tag_949.re;
  assign rcache_line[3][181].status_reg.status = reg2hw.status_949.q;//status_reg_t'(reg2hw.status_949.q);
  assign rcache_line[3][181].status_reg.qe    = reg2hw.status_949.qe;
  assign rcache_line[3][181].status_reg.re    = reg2hw.status_949.re;


  assign rcache_line[3][182].tag_reg.tag      = reg2hw.tag_950.q;
  assign rcache_line[3][182].tag_reg.qe       = reg2hw.tag_950.qe;
  assign rcache_line[3][182].tag_reg.re       = reg2hw.tag_950.re;
  assign rcache_line[3][182].status_reg.status = reg2hw.status_950.q;//status_reg_t'(reg2hw.status_950.q);
  assign rcache_line[3][182].status_reg.qe    = reg2hw.status_950.qe;
  assign rcache_line[3][182].status_reg.re    = reg2hw.status_950.re;


  assign rcache_line[3][183].tag_reg.tag      = reg2hw.tag_951.q;
  assign rcache_line[3][183].tag_reg.qe       = reg2hw.tag_951.qe;
  assign rcache_line[3][183].tag_reg.re       = reg2hw.tag_951.re;
  assign rcache_line[3][183].status_reg.status = reg2hw.status_951.q;//status_reg_t'(reg2hw.status_951.q);
  assign rcache_line[3][183].status_reg.qe    = reg2hw.status_951.qe;
  assign rcache_line[3][183].status_reg.re    = reg2hw.status_951.re;


  assign rcache_line[3][184].tag_reg.tag      = reg2hw.tag_952.q;
  assign rcache_line[3][184].tag_reg.qe       = reg2hw.tag_952.qe;
  assign rcache_line[3][184].tag_reg.re       = reg2hw.tag_952.re;
  assign rcache_line[3][184].status_reg.status = reg2hw.status_952.q;//status_reg_t'(reg2hw.status_952.q);
  assign rcache_line[3][184].status_reg.qe    = reg2hw.status_952.qe;
  assign rcache_line[3][184].status_reg.re    = reg2hw.status_952.re;


  assign rcache_line[3][185].tag_reg.tag      = reg2hw.tag_953.q;
  assign rcache_line[3][185].tag_reg.qe       = reg2hw.tag_953.qe;
  assign rcache_line[3][185].tag_reg.re       = reg2hw.tag_953.re;
  assign rcache_line[3][185].status_reg.status = reg2hw.status_953.q;//status_reg_t'(reg2hw.status_953.q);
  assign rcache_line[3][185].status_reg.qe    = reg2hw.status_953.qe;
  assign rcache_line[3][185].status_reg.re    = reg2hw.status_953.re;


  assign rcache_line[3][186].tag_reg.tag      = reg2hw.tag_954.q;
  assign rcache_line[3][186].tag_reg.qe       = reg2hw.tag_954.qe;
  assign rcache_line[3][186].tag_reg.re       = reg2hw.tag_954.re;
  assign rcache_line[3][186].status_reg.status = reg2hw.status_954.q;//status_reg_t'(reg2hw.status_954.q);
  assign rcache_line[3][186].status_reg.qe    = reg2hw.status_954.qe;
  assign rcache_line[3][186].status_reg.re    = reg2hw.status_954.re;


  assign rcache_line[3][187].tag_reg.tag      = reg2hw.tag_955.q;
  assign rcache_line[3][187].tag_reg.qe       = reg2hw.tag_955.qe;
  assign rcache_line[3][187].tag_reg.re       = reg2hw.tag_955.re;
  assign rcache_line[3][187].status_reg.status = reg2hw.status_955.q;//status_reg_t'(reg2hw.status_955.q);
  assign rcache_line[3][187].status_reg.qe    = reg2hw.status_955.qe;
  assign rcache_line[3][187].status_reg.re    = reg2hw.status_955.re;


  assign rcache_line[3][188].tag_reg.tag      = reg2hw.tag_956.q;
  assign rcache_line[3][188].tag_reg.qe       = reg2hw.tag_956.qe;
  assign rcache_line[3][188].tag_reg.re       = reg2hw.tag_956.re;
  assign rcache_line[3][188].status_reg.status = reg2hw.status_956.q;//status_reg_t'(reg2hw.status_956.q);
  assign rcache_line[3][188].status_reg.qe    = reg2hw.status_956.qe;
  assign rcache_line[3][188].status_reg.re    = reg2hw.status_956.re;


  assign rcache_line[3][189].tag_reg.tag      = reg2hw.tag_957.q;
  assign rcache_line[3][189].tag_reg.qe       = reg2hw.tag_957.qe;
  assign rcache_line[3][189].tag_reg.re       = reg2hw.tag_957.re;
  assign rcache_line[3][189].status_reg.status = reg2hw.status_957.q;//status_reg_t'(reg2hw.status_957.q);
  assign rcache_line[3][189].status_reg.qe    = reg2hw.status_957.qe;
  assign rcache_line[3][189].status_reg.re    = reg2hw.status_957.re;


  assign rcache_line[3][190].tag_reg.tag      = reg2hw.tag_958.q;
  assign rcache_line[3][190].tag_reg.qe       = reg2hw.tag_958.qe;
  assign rcache_line[3][190].tag_reg.re       = reg2hw.tag_958.re;
  assign rcache_line[3][190].status_reg.status = reg2hw.status_958.q;//status_reg_t'(reg2hw.status_958.q);
  assign rcache_line[3][190].status_reg.qe    = reg2hw.status_958.qe;
  assign rcache_line[3][190].status_reg.re    = reg2hw.status_958.re;


  assign rcache_line[3][191].tag_reg.tag      = reg2hw.tag_959.q;
  assign rcache_line[3][191].tag_reg.qe       = reg2hw.tag_959.qe;
  assign rcache_line[3][191].tag_reg.re       = reg2hw.tag_959.re;
  assign rcache_line[3][191].status_reg.status = reg2hw.status_959.q;//status_reg_t'(reg2hw.status_959.q);
  assign rcache_line[3][191].status_reg.qe    = reg2hw.status_959.qe;
  assign rcache_line[3][191].status_reg.re    = reg2hw.status_959.re;


  assign rcache_line[3][192].tag_reg.tag      = reg2hw.tag_960.q;
  assign rcache_line[3][192].tag_reg.qe       = reg2hw.tag_960.qe;
  assign rcache_line[3][192].tag_reg.re       = reg2hw.tag_960.re;
  assign rcache_line[3][192].status_reg.status = reg2hw.status_960.q;//status_reg_t'(reg2hw.status_960.q);
  assign rcache_line[3][192].status_reg.qe    = reg2hw.status_960.qe;
  assign rcache_line[3][192].status_reg.re    = reg2hw.status_960.re;


  assign rcache_line[3][193].tag_reg.tag      = reg2hw.tag_961.q;
  assign rcache_line[3][193].tag_reg.qe       = reg2hw.tag_961.qe;
  assign rcache_line[3][193].tag_reg.re       = reg2hw.tag_961.re;
  assign rcache_line[3][193].status_reg.status = reg2hw.status_961.q;//status_reg_t'(reg2hw.status_961.q);
  assign rcache_line[3][193].status_reg.qe    = reg2hw.status_961.qe;
  assign rcache_line[3][193].status_reg.re    = reg2hw.status_961.re;


  assign rcache_line[3][194].tag_reg.tag      = reg2hw.tag_962.q;
  assign rcache_line[3][194].tag_reg.qe       = reg2hw.tag_962.qe;
  assign rcache_line[3][194].tag_reg.re       = reg2hw.tag_962.re;
  assign rcache_line[3][194].status_reg.status = reg2hw.status_962.q;//status_reg_t'(reg2hw.status_962.q);
  assign rcache_line[3][194].status_reg.qe    = reg2hw.status_962.qe;
  assign rcache_line[3][194].status_reg.re    = reg2hw.status_962.re;


  assign rcache_line[3][195].tag_reg.tag      = reg2hw.tag_963.q;
  assign rcache_line[3][195].tag_reg.qe       = reg2hw.tag_963.qe;
  assign rcache_line[3][195].tag_reg.re       = reg2hw.tag_963.re;
  assign rcache_line[3][195].status_reg.status = reg2hw.status_963.q;//status_reg_t'(reg2hw.status_963.q);
  assign rcache_line[3][195].status_reg.qe    = reg2hw.status_963.qe;
  assign rcache_line[3][195].status_reg.re    = reg2hw.status_963.re;


  assign rcache_line[3][196].tag_reg.tag      = reg2hw.tag_964.q;
  assign rcache_line[3][196].tag_reg.qe       = reg2hw.tag_964.qe;
  assign rcache_line[3][196].tag_reg.re       = reg2hw.tag_964.re;
  assign rcache_line[3][196].status_reg.status = reg2hw.status_964.q;//status_reg_t'(reg2hw.status_964.q);
  assign rcache_line[3][196].status_reg.qe    = reg2hw.status_964.qe;
  assign rcache_line[3][196].status_reg.re    = reg2hw.status_964.re;


  assign rcache_line[3][197].tag_reg.tag      = reg2hw.tag_965.q;
  assign rcache_line[3][197].tag_reg.qe       = reg2hw.tag_965.qe;
  assign rcache_line[3][197].tag_reg.re       = reg2hw.tag_965.re;
  assign rcache_line[3][197].status_reg.status = reg2hw.status_965.q;//status_reg_t'(reg2hw.status_965.q);
  assign rcache_line[3][197].status_reg.qe    = reg2hw.status_965.qe;
  assign rcache_line[3][197].status_reg.re    = reg2hw.status_965.re;


  assign rcache_line[3][198].tag_reg.tag      = reg2hw.tag_966.q;
  assign rcache_line[3][198].tag_reg.qe       = reg2hw.tag_966.qe;
  assign rcache_line[3][198].tag_reg.re       = reg2hw.tag_966.re;
  assign rcache_line[3][198].status_reg.status = reg2hw.status_966.q;//status_reg_t'(reg2hw.status_966.q);
  assign rcache_line[3][198].status_reg.qe    = reg2hw.status_966.qe;
  assign rcache_line[3][198].status_reg.re    = reg2hw.status_966.re;


  assign rcache_line[3][199].tag_reg.tag      = reg2hw.tag_967.q;
  assign rcache_line[3][199].tag_reg.qe       = reg2hw.tag_967.qe;
  assign rcache_line[3][199].tag_reg.re       = reg2hw.tag_967.re;
  assign rcache_line[3][199].status_reg.status = reg2hw.status_967.q;//status_reg_t'(reg2hw.status_967.q);
  assign rcache_line[3][199].status_reg.qe    = reg2hw.status_967.qe;
  assign rcache_line[3][199].status_reg.re    = reg2hw.status_967.re;


  assign rcache_line[3][200].tag_reg.tag      = reg2hw.tag_968.q;
  assign rcache_line[3][200].tag_reg.qe       = reg2hw.tag_968.qe;
  assign rcache_line[3][200].tag_reg.re       = reg2hw.tag_968.re;
  assign rcache_line[3][200].status_reg.status = reg2hw.status_968.q;//status_reg_t'(reg2hw.status_968.q);
  assign rcache_line[3][200].status_reg.qe    = reg2hw.status_968.qe;
  assign rcache_line[3][200].status_reg.re    = reg2hw.status_968.re;


  assign rcache_line[3][201].tag_reg.tag      = reg2hw.tag_969.q;
  assign rcache_line[3][201].tag_reg.qe       = reg2hw.tag_969.qe;
  assign rcache_line[3][201].tag_reg.re       = reg2hw.tag_969.re;
  assign rcache_line[3][201].status_reg.status = reg2hw.status_969.q;//status_reg_t'(reg2hw.status_969.q);
  assign rcache_line[3][201].status_reg.qe    = reg2hw.status_969.qe;
  assign rcache_line[3][201].status_reg.re    = reg2hw.status_969.re;


  assign rcache_line[3][202].tag_reg.tag      = reg2hw.tag_970.q;
  assign rcache_line[3][202].tag_reg.qe       = reg2hw.tag_970.qe;
  assign rcache_line[3][202].tag_reg.re       = reg2hw.tag_970.re;
  assign rcache_line[3][202].status_reg.status = reg2hw.status_970.q;//status_reg_t'(reg2hw.status_970.q);
  assign rcache_line[3][202].status_reg.qe    = reg2hw.status_970.qe;
  assign rcache_line[3][202].status_reg.re    = reg2hw.status_970.re;


  assign rcache_line[3][203].tag_reg.tag      = reg2hw.tag_971.q;
  assign rcache_line[3][203].tag_reg.qe       = reg2hw.tag_971.qe;
  assign rcache_line[3][203].tag_reg.re       = reg2hw.tag_971.re;
  assign rcache_line[3][203].status_reg.status = reg2hw.status_971.q;//status_reg_t'(reg2hw.status_971.q);
  assign rcache_line[3][203].status_reg.qe    = reg2hw.status_971.qe;
  assign rcache_line[3][203].status_reg.re    = reg2hw.status_971.re;


  assign rcache_line[3][204].tag_reg.tag      = reg2hw.tag_972.q;
  assign rcache_line[3][204].tag_reg.qe       = reg2hw.tag_972.qe;
  assign rcache_line[3][204].tag_reg.re       = reg2hw.tag_972.re;
  assign rcache_line[3][204].status_reg.status = reg2hw.status_972.q;//status_reg_t'(reg2hw.status_972.q);
  assign rcache_line[3][204].status_reg.qe    = reg2hw.status_972.qe;
  assign rcache_line[3][204].status_reg.re    = reg2hw.status_972.re;


  assign rcache_line[3][205].tag_reg.tag      = reg2hw.tag_973.q;
  assign rcache_line[3][205].tag_reg.qe       = reg2hw.tag_973.qe;
  assign rcache_line[3][205].tag_reg.re       = reg2hw.tag_973.re;
  assign rcache_line[3][205].status_reg.status = reg2hw.status_973.q;//status_reg_t'(reg2hw.status_973.q);
  assign rcache_line[3][205].status_reg.qe    = reg2hw.status_973.qe;
  assign rcache_line[3][205].status_reg.re    = reg2hw.status_973.re;


  assign rcache_line[3][206].tag_reg.tag      = reg2hw.tag_974.q;
  assign rcache_line[3][206].tag_reg.qe       = reg2hw.tag_974.qe;
  assign rcache_line[3][206].tag_reg.re       = reg2hw.tag_974.re;
  assign rcache_line[3][206].status_reg.status = reg2hw.status_974.q;//status_reg_t'(reg2hw.status_974.q);
  assign rcache_line[3][206].status_reg.qe    = reg2hw.status_974.qe;
  assign rcache_line[3][206].status_reg.re    = reg2hw.status_974.re;


  assign rcache_line[3][207].tag_reg.tag      = reg2hw.tag_975.q;
  assign rcache_line[3][207].tag_reg.qe       = reg2hw.tag_975.qe;
  assign rcache_line[3][207].tag_reg.re       = reg2hw.tag_975.re;
  assign rcache_line[3][207].status_reg.status = reg2hw.status_975.q;//status_reg_t'(reg2hw.status_975.q);
  assign rcache_line[3][207].status_reg.qe    = reg2hw.status_975.qe;
  assign rcache_line[3][207].status_reg.re    = reg2hw.status_975.re;


  assign rcache_line[3][208].tag_reg.tag      = reg2hw.tag_976.q;
  assign rcache_line[3][208].tag_reg.qe       = reg2hw.tag_976.qe;
  assign rcache_line[3][208].tag_reg.re       = reg2hw.tag_976.re;
  assign rcache_line[3][208].status_reg.status = reg2hw.status_976.q;//status_reg_t'(reg2hw.status_976.q);
  assign rcache_line[3][208].status_reg.qe    = reg2hw.status_976.qe;
  assign rcache_line[3][208].status_reg.re    = reg2hw.status_976.re;


  assign rcache_line[3][209].tag_reg.tag      = reg2hw.tag_977.q;
  assign rcache_line[3][209].tag_reg.qe       = reg2hw.tag_977.qe;
  assign rcache_line[3][209].tag_reg.re       = reg2hw.tag_977.re;
  assign rcache_line[3][209].status_reg.status = reg2hw.status_977.q;//status_reg_t'(reg2hw.status_977.q);
  assign rcache_line[3][209].status_reg.qe    = reg2hw.status_977.qe;
  assign rcache_line[3][209].status_reg.re    = reg2hw.status_977.re;


  assign rcache_line[3][210].tag_reg.tag      = reg2hw.tag_978.q;
  assign rcache_line[3][210].tag_reg.qe       = reg2hw.tag_978.qe;
  assign rcache_line[3][210].tag_reg.re       = reg2hw.tag_978.re;
  assign rcache_line[3][210].status_reg.status = reg2hw.status_978.q;//status_reg_t'(reg2hw.status_978.q);
  assign rcache_line[3][210].status_reg.qe    = reg2hw.status_978.qe;
  assign rcache_line[3][210].status_reg.re    = reg2hw.status_978.re;


  assign rcache_line[3][211].tag_reg.tag      = reg2hw.tag_979.q;
  assign rcache_line[3][211].tag_reg.qe       = reg2hw.tag_979.qe;
  assign rcache_line[3][211].tag_reg.re       = reg2hw.tag_979.re;
  assign rcache_line[3][211].status_reg.status = reg2hw.status_979.q;//status_reg_t'(reg2hw.status_979.q);
  assign rcache_line[3][211].status_reg.qe    = reg2hw.status_979.qe;
  assign rcache_line[3][211].status_reg.re    = reg2hw.status_979.re;


  assign rcache_line[3][212].tag_reg.tag      = reg2hw.tag_980.q;
  assign rcache_line[3][212].tag_reg.qe       = reg2hw.tag_980.qe;
  assign rcache_line[3][212].tag_reg.re       = reg2hw.tag_980.re;
  assign rcache_line[3][212].status_reg.status = reg2hw.status_980.q;//status_reg_t'(reg2hw.status_980.q);
  assign rcache_line[3][212].status_reg.qe    = reg2hw.status_980.qe;
  assign rcache_line[3][212].status_reg.re    = reg2hw.status_980.re;


  assign rcache_line[3][213].tag_reg.tag      = reg2hw.tag_981.q;
  assign rcache_line[3][213].tag_reg.qe       = reg2hw.tag_981.qe;
  assign rcache_line[3][213].tag_reg.re       = reg2hw.tag_981.re;
  assign rcache_line[3][213].status_reg.status = reg2hw.status_981.q;//status_reg_t'(reg2hw.status_981.q);
  assign rcache_line[3][213].status_reg.qe    = reg2hw.status_981.qe;
  assign rcache_line[3][213].status_reg.re    = reg2hw.status_981.re;


  assign rcache_line[3][214].tag_reg.tag      = reg2hw.tag_982.q;
  assign rcache_line[3][214].tag_reg.qe       = reg2hw.tag_982.qe;
  assign rcache_line[3][214].tag_reg.re       = reg2hw.tag_982.re;
  assign rcache_line[3][214].status_reg.status = reg2hw.status_982.q;//status_reg_t'(reg2hw.status_982.q);
  assign rcache_line[3][214].status_reg.qe    = reg2hw.status_982.qe;
  assign rcache_line[3][214].status_reg.re    = reg2hw.status_982.re;


  assign rcache_line[3][215].tag_reg.tag      = reg2hw.tag_983.q;
  assign rcache_line[3][215].tag_reg.qe       = reg2hw.tag_983.qe;
  assign rcache_line[3][215].tag_reg.re       = reg2hw.tag_983.re;
  assign rcache_line[3][215].status_reg.status = reg2hw.status_983.q;//status_reg_t'(reg2hw.status_983.q);
  assign rcache_line[3][215].status_reg.qe    = reg2hw.status_983.qe;
  assign rcache_line[3][215].status_reg.re    = reg2hw.status_983.re;


  assign rcache_line[3][216].tag_reg.tag      = reg2hw.tag_984.q;
  assign rcache_line[3][216].tag_reg.qe       = reg2hw.tag_984.qe;
  assign rcache_line[3][216].tag_reg.re       = reg2hw.tag_984.re;
  assign rcache_line[3][216].status_reg.status = reg2hw.status_984.q;//status_reg_t'(reg2hw.status_984.q);
  assign rcache_line[3][216].status_reg.qe    = reg2hw.status_984.qe;
  assign rcache_line[3][216].status_reg.re    = reg2hw.status_984.re;


  assign rcache_line[3][217].tag_reg.tag      = reg2hw.tag_985.q;
  assign rcache_line[3][217].tag_reg.qe       = reg2hw.tag_985.qe;
  assign rcache_line[3][217].tag_reg.re       = reg2hw.tag_985.re;
  assign rcache_line[3][217].status_reg.status = reg2hw.status_985.q;//status_reg_t'(reg2hw.status_985.q);
  assign rcache_line[3][217].status_reg.qe    = reg2hw.status_985.qe;
  assign rcache_line[3][217].status_reg.re    = reg2hw.status_985.re;


  assign rcache_line[3][218].tag_reg.tag      = reg2hw.tag_986.q;
  assign rcache_line[3][218].tag_reg.qe       = reg2hw.tag_986.qe;
  assign rcache_line[3][218].tag_reg.re       = reg2hw.tag_986.re;
  assign rcache_line[3][218].status_reg.status = reg2hw.status_986.q;//status_reg_t'(reg2hw.status_986.q);
  assign rcache_line[3][218].status_reg.qe    = reg2hw.status_986.qe;
  assign rcache_line[3][218].status_reg.re    = reg2hw.status_986.re;


  assign rcache_line[3][219].tag_reg.tag      = reg2hw.tag_987.q;
  assign rcache_line[3][219].tag_reg.qe       = reg2hw.tag_987.qe;
  assign rcache_line[3][219].tag_reg.re       = reg2hw.tag_987.re;
  assign rcache_line[3][219].status_reg.status = reg2hw.status_987.q;//status_reg_t'(reg2hw.status_987.q);
  assign rcache_line[3][219].status_reg.qe    = reg2hw.status_987.qe;
  assign rcache_line[3][219].status_reg.re    = reg2hw.status_987.re;


  assign rcache_line[3][220].tag_reg.tag      = reg2hw.tag_988.q;
  assign rcache_line[3][220].tag_reg.qe       = reg2hw.tag_988.qe;
  assign rcache_line[3][220].tag_reg.re       = reg2hw.tag_988.re;
  assign rcache_line[3][220].status_reg.status = reg2hw.status_988.q;//status_reg_t'(reg2hw.status_988.q);
  assign rcache_line[3][220].status_reg.qe    = reg2hw.status_988.qe;
  assign rcache_line[3][220].status_reg.re    = reg2hw.status_988.re;


  assign rcache_line[3][221].tag_reg.tag      = reg2hw.tag_989.q;
  assign rcache_line[3][221].tag_reg.qe       = reg2hw.tag_989.qe;
  assign rcache_line[3][221].tag_reg.re       = reg2hw.tag_989.re;
  assign rcache_line[3][221].status_reg.status = reg2hw.status_989.q;//status_reg_t'(reg2hw.status_989.q);
  assign rcache_line[3][221].status_reg.qe    = reg2hw.status_989.qe;
  assign rcache_line[3][221].status_reg.re    = reg2hw.status_989.re;


  assign rcache_line[3][222].tag_reg.tag      = reg2hw.tag_990.q;
  assign rcache_line[3][222].tag_reg.qe       = reg2hw.tag_990.qe;
  assign rcache_line[3][222].tag_reg.re       = reg2hw.tag_990.re;
  assign rcache_line[3][222].status_reg.status = reg2hw.status_990.q;//status_reg_t'(reg2hw.status_990.q);
  assign rcache_line[3][222].status_reg.qe    = reg2hw.status_990.qe;
  assign rcache_line[3][222].status_reg.re    = reg2hw.status_990.re;


  assign rcache_line[3][223].tag_reg.tag      = reg2hw.tag_991.q;
  assign rcache_line[3][223].tag_reg.qe       = reg2hw.tag_991.qe;
  assign rcache_line[3][223].tag_reg.re       = reg2hw.tag_991.re;
  assign rcache_line[3][223].status_reg.status = reg2hw.status_991.q;//status_reg_t'(reg2hw.status_991.q);
  assign rcache_line[3][223].status_reg.qe    = reg2hw.status_991.qe;
  assign rcache_line[3][223].status_reg.re    = reg2hw.status_991.re;


  assign rcache_line[3][224].tag_reg.tag      = reg2hw.tag_992.q;
  assign rcache_line[3][224].tag_reg.qe       = reg2hw.tag_992.qe;
  assign rcache_line[3][224].tag_reg.re       = reg2hw.tag_992.re;
  assign rcache_line[3][224].status_reg.status = reg2hw.status_992.q;//status_reg_t'(reg2hw.status_992.q);
  assign rcache_line[3][224].status_reg.qe    = reg2hw.status_992.qe;
  assign rcache_line[3][224].status_reg.re    = reg2hw.status_992.re;


  assign rcache_line[3][225].tag_reg.tag      = reg2hw.tag_993.q;
  assign rcache_line[3][225].tag_reg.qe       = reg2hw.tag_993.qe;
  assign rcache_line[3][225].tag_reg.re       = reg2hw.tag_993.re;
  assign rcache_line[3][225].status_reg.status = reg2hw.status_993.q;//status_reg_t'(reg2hw.status_993.q);
  assign rcache_line[3][225].status_reg.qe    = reg2hw.status_993.qe;
  assign rcache_line[3][225].status_reg.re    = reg2hw.status_993.re;


  assign rcache_line[3][226].tag_reg.tag      = reg2hw.tag_994.q;
  assign rcache_line[3][226].tag_reg.qe       = reg2hw.tag_994.qe;
  assign rcache_line[3][226].tag_reg.re       = reg2hw.tag_994.re;
  assign rcache_line[3][226].status_reg.status = reg2hw.status_994.q;//status_reg_t'(reg2hw.status_994.q);
  assign rcache_line[3][226].status_reg.qe    = reg2hw.status_994.qe;
  assign rcache_line[3][226].status_reg.re    = reg2hw.status_994.re;


  assign rcache_line[3][227].tag_reg.tag      = reg2hw.tag_995.q;
  assign rcache_line[3][227].tag_reg.qe       = reg2hw.tag_995.qe;
  assign rcache_line[3][227].tag_reg.re       = reg2hw.tag_995.re;
  assign rcache_line[3][227].status_reg.status = reg2hw.status_995.q;//status_reg_t'(reg2hw.status_995.q);
  assign rcache_line[3][227].status_reg.qe    = reg2hw.status_995.qe;
  assign rcache_line[3][227].status_reg.re    = reg2hw.status_995.re;


  assign rcache_line[3][228].tag_reg.tag      = reg2hw.tag_996.q;
  assign rcache_line[3][228].tag_reg.qe       = reg2hw.tag_996.qe;
  assign rcache_line[3][228].tag_reg.re       = reg2hw.tag_996.re;
  assign rcache_line[3][228].status_reg.status = reg2hw.status_996.q;//status_reg_t'(reg2hw.status_996.q);
  assign rcache_line[3][228].status_reg.qe    = reg2hw.status_996.qe;
  assign rcache_line[3][228].status_reg.re    = reg2hw.status_996.re;


  assign rcache_line[3][229].tag_reg.tag      = reg2hw.tag_997.q;
  assign rcache_line[3][229].tag_reg.qe       = reg2hw.tag_997.qe;
  assign rcache_line[3][229].tag_reg.re       = reg2hw.tag_997.re;
  assign rcache_line[3][229].status_reg.status = reg2hw.status_997.q;//status_reg_t'(reg2hw.status_997.q);
  assign rcache_line[3][229].status_reg.qe    = reg2hw.status_997.qe;
  assign rcache_line[3][229].status_reg.re    = reg2hw.status_997.re;


  assign rcache_line[3][230].tag_reg.tag      = reg2hw.tag_998.q;
  assign rcache_line[3][230].tag_reg.qe       = reg2hw.tag_998.qe;
  assign rcache_line[3][230].tag_reg.re       = reg2hw.tag_998.re;
  assign rcache_line[3][230].status_reg.status = reg2hw.status_998.q;//status_reg_t'(reg2hw.status_998.q);
  assign rcache_line[3][230].status_reg.qe    = reg2hw.status_998.qe;
  assign rcache_line[3][230].status_reg.re    = reg2hw.status_998.re;


  assign rcache_line[3][231].tag_reg.tag      = reg2hw.tag_999.q;
  assign rcache_line[3][231].tag_reg.qe       = reg2hw.tag_999.qe;
  assign rcache_line[3][231].tag_reg.re       = reg2hw.tag_999.re;
  assign rcache_line[3][231].status_reg.status = reg2hw.status_999.q;//status_reg_t'(reg2hw.status_999.q);
  assign rcache_line[3][231].status_reg.qe    = reg2hw.status_999.qe;
  assign rcache_line[3][231].status_reg.re    = reg2hw.status_999.re;


  assign rcache_line[3][232].tag_reg.tag      = reg2hw.tag_1000.q;
  assign rcache_line[3][232].tag_reg.qe       = reg2hw.tag_1000.qe;
  assign rcache_line[3][232].tag_reg.re       = reg2hw.tag_1000.re;
  assign rcache_line[3][232].status_reg.status = reg2hw.status_1000.q;//status_reg_t'(reg2hw.status_1000.q);
  assign rcache_line[3][232].status_reg.qe    = reg2hw.status_1000.qe;
  assign rcache_line[3][232].status_reg.re    = reg2hw.status_1000.re;


  assign rcache_line[3][233].tag_reg.tag      = reg2hw.tag_1001.q;
  assign rcache_line[3][233].tag_reg.qe       = reg2hw.tag_1001.qe;
  assign rcache_line[3][233].tag_reg.re       = reg2hw.tag_1001.re;
  assign rcache_line[3][233].status_reg.status = reg2hw.status_1001.q;//status_reg_t'(reg2hw.status_1001.q);
  assign rcache_line[3][233].status_reg.qe    = reg2hw.status_1001.qe;
  assign rcache_line[3][233].status_reg.re    = reg2hw.status_1001.re;


  assign rcache_line[3][234].tag_reg.tag      = reg2hw.tag_1002.q;
  assign rcache_line[3][234].tag_reg.qe       = reg2hw.tag_1002.qe;
  assign rcache_line[3][234].tag_reg.re       = reg2hw.tag_1002.re;
  assign rcache_line[3][234].status_reg.status = reg2hw.status_1002.q;//status_reg_t'(reg2hw.status_1002.q);
  assign rcache_line[3][234].status_reg.qe    = reg2hw.status_1002.qe;
  assign rcache_line[3][234].status_reg.re    = reg2hw.status_1002.re;


  assign rcache_line[3][235].tag_reg.tag      = reg2hw.tag_1003.q;
  assign rcache_line[3][235].tag_reg.qe       = reg2hw.tag_1003.qe;
  assign rcache_line[3][235].tag_reg.re       = reg2hw.tag_1003.re;
  assign rcache_line[3][235].status_reg.status = reg2hw.status_1003.q;//status_reg_t'(reg2hw.status_1003.q);
  assign rcache_line[3][235].status_reg.qe    = reg2hw.status_1003.qe;
  assign rcache_line[3][235].status_reg.re    = reg2hw.status_1003.re;


  assign rcache_line[3][236].tag_reg.tag      = reg2hw.tag_1004.q;
  assign rcache_line[3][236].tag_reg.qe       = reg2hw.tag_1004.qe;
  assign rcache_line[3][236].tag_reg.re       = reg2hw.tag_1004.re;
  assign rcache_line[3][236].status_reg.status = reg2hw.status_1004.q;//status_reg_t'(reg2hw.status_1004.q);
  assign rcache_line[3][236].status_reg.qe    = reg2hw.status_1004.qe;
  assign rcache_line[3][236].status_reg.re    = reg2hw.status_1004.re;


  assign rcache_line[3][237].tag_reg.tag      = reg2hw.tag_1005.q;
  assign rcache_line[3][237].tag_reg.qe       = reg2hw.tag_1005.qe;
  assign rcache_line[3][237].tag_reg.re       = reg2hw.tag_1005.re;
  assign rcache_line[3][237].status_reg.status = reg2hw.status_1005.q;//status_reg_t'(reg2hw.status_1005.q);
  assign rcache_line[3][237].status_reg.qe    = reg2hw.status_1005.qe;
  assign rcache_line[3][237].status_reg.re    = reg2hw.status_1005.re;


  assign rcache_line[3][238].tag_reg.tag      = reg2hw.tag_1006.q;
  assign rcache_line[3][238].tag_reg.qe       = reg2hw.tag_1006.qe;
  assign rcache_line[3][238].tag_reg.re       = reg2hw.tag_1006.re;
  assign rcache_line[3][238].status_reg.status = reg2hw.status_1006.q;//status_reg_t'(reg2hw.status_1006.q);
  assign rcache_line[3][238].status_reg.qe    = reg2hw.status_1006.qe;
  assign rcache_line[3][238].status_reg.re    = reg2hw.status_1006.re;


  assign rcache_line[3][239].tag_reg.tag      = reg2hw.tag_1007.q;
  assign rcache_line[3][239].tag_reg.qe       = reg2hw.tag_1007.qe;
  assign rcache_line[3][239].tag_reg.re       = reg2hw.tag_1007.re;
  assign rcache_line[3][239].status_reg.status = reg2hw.status_1007.q;//status_reg_t'(reg2hw.status_1007.q);
  assign rcache_line[3][239].status_reg.qe    = reg2hw.status_1007.qe;
  assign rcache_line[3][239].status_reg.re    = reg2hw.status_1007.re;


  assign rcache_line[3][240].tag_reg.tag      = reg2hw.tag_1008.q;
  assign rcache_line[3][240].tag_reg.qe       = reg2hw.tag_1008.qe;
  assign rcache_line[3][240].tag_reg.re       = reg2hw.tag_1008.re;
  assign rcache_line[3][240].status_reg.status = reg2hw.status_1008.q;//status_reg_t'(reg2hw.status_1008.q);
  assign rcache_line[3][240].status_reg.qe    = reg2hw.status_1008.qe;
  assign rcache_line[3][240].status_reg.re    = reg2hw.status_1008.re;


  assign rcache_line[3][241].tag_reg.tag      = reg2hw.tag_1009.q;
  assign rcache_line[3][241].tag_reg.qe       = reg2hw.tag_1009.qe;
  assign rcache_line[3][241].tag_reg.re       = reg2hw.tag_1009.re;
  assign rcache_line[3][241].status_reg.status = reg2hw.status_1009.q;//status_reg_t'(reg2hw.status_1009.q);
  assign rcache_line[3][241].status_reg.qe    = reg2hw.status_1009.qe;
  assign rcache_line[3][241].status_reg.re    = reg2hw.status_1009.re;


  assign rcache_line[3][242].tag_reg.tag      = reg2hw.tag_1010.q;
  assign rcache_line[3][242].tag_reg.qe       = reg2hw.tag_1010.qe;
  assign rcache_line[3][242].tag_reg.re       = reg2hw.tag_1010.re;
  assign rcache_line[3][242].status_reg.status = reg2hw.status_1010.q;//status_reg_t'(reg2hw.status_1010.q);
  assign rcache_line[3][242].status_reg.qe    = reg2hw.status_1010.qe;
  assign rcache_line[3][242].status_reg.re    = reg2hw.status_1010.re;


  assign rcache_line[3][243].tag_reg.tag      = reg2hw.tag_1011.q;
  assign rcache_line[3][243].tag_reg.qe       = reg2hw.tag_1011.qe;
  assign rcache_line[3][243].tag_reg.re       = reg2hw.tag_1011.re;
  assign rcache_line[3][243].status_reg.status = reg2hw.status_1011.q;//status_reg_t'(reg2hw.status_1011.q);
  assign rcache_line[3][243].status_reg.qe    = reg2hw.status_1011.qe;
  assign rcache_line[3][243].status_reg.re    = reg2hw.status_1011.re;


  assign rcache_line[3][244].tag_reg.tag      = reg2hw.tag_1012.q;
  assign rcache_line[3][244].tag_reg.qe       = reg2hw.tag_1012.qe;
  assign rcache_line[3][244].tag_reg.re       = reg2hw.tag_1012.re;
  assign rcache_line[3][244].status_reg.status = reg2hw.status_1012.q;//status_reg_t'(reg2hw.status_1012.q);
  assign rcache_line[3][244].status_reg.qe    = reg2hw.status_1012.qe;
  assign rcache_line[3][244].status_reg.re    = reg2hw.status_1012.re;


  assign rcache_line[3][245].tag_reg.tag      = reg2hw.tag_1013.q;
  assign rcache_line[3][245].tag_reg.qe       = reg2hw.tag_1013.qe;
  assign rcache_line[3][245].tag_reg.re       = reg2hw.tag_1013.re;
  assign rcache_line[3][245].status_reg.status = reg2hw.status_1013.q;//status_reg_t'(reg2hw.status_1013.q);
  assign rcache_line[3][245].status_reg.qe    = reg2hw.status_1013.qe;
  assign rcache_line[3][245].status_reg.re    = reg2hw.status_1013.re;


  assign rcache_line[3][246].tag_reg.tag      = reg2hw.tag_1014.q;
  assign rcache_line[3][246].tag_reg.qe       = reg2hw.tag_1014.qe;
  assign rcache_line[3][246].tag_reg.re       = reg2hw.tag_1014.re;
  assign rcache_line[3][246].status_reg.status = reg2hw.status_1014.q;//status_reg_t'(reg2hw.status_1014.q);
  assign rcache_line[3][246].status_reg.qe    = reg2hw.status_1014.qe;
  assign rcache_line[3][246].status_reg.re    = reg2hw.status_1014.re;


  assign rcache_line[3][247].tag_reg.tag      = reg2hw.tag_1015.q;
  assign rcache_line[3][247].tag_reg.qe       = reg2hw.tag_1015.qe;
  assign rcache_line[3][247].tag_reg.re       = reg2hw.tag_1015.re;
  assign rcache_line[3][247].status_reg.status = reg2hw.status_1015.q;//status_reg_t'(reg2hw.status_1015.q);
  assign rcache_line[3][247].status_reg.qe    = reg2hw.status_1015.qe;
  assign rcache_line[3][247].status_reg.re    = reg2hw.status_1015.re;


  assign rcache_line[3][248].tag_reg.tag      = reg2hw.tag_1016.q;
  assign rcache_line[3][248].tag_reg.qe       = reg2hw.tag_1016.qe;
  assign rcache_line[3][248].tag_reg.re       = reg2hw.tag_1016.re;
  assign rcache_line[3][248].status_reg.status = reg2hw.status_1016.q;//status_reg_t'(reg2hw.status_1016.q);
  assign rcache_line[3][248].status_reg.qe    = reg2hw.status_1016.qe;
  assign rcache_line[3][248].status_reg.re    = reg2hw.status_1016.re;


  assign rcache_line[3][249].tag_reg.tag      = reg2hw.tag_1017.q;
  assign rcache_line[3][249].tag_reg.qe       = reg2hw.tag_1017.qe;
  assign rcache_line[3][249].tag_reg.re       = reg2hw.tag_1017.re;
  assign rcache_line[3][249].status_reg.status = reg2hw.status_1017.q;//status_reg_t'(reg2hw.status_1017.q);
  assign rcache_line[3][249].status_reg.qe    = reg2hw.status_1017.qe;
  assign rcache_line[3][249].status_reg.re    = reg2hw.status_1017.re;


  assign rcache_line[3][250].tag_reg.tag      = reg2hw.tag_1018.q;
  assign rcache_line[3][250].tag_reg.qe       = reg2hw.tag_1018.qe;
  assign rcache_line[3][250].tag_reg.re       = reg2hw.tag_1018.re;
  assign rcache_line[3][250].status_reg.status = reg2hw.status_1018.q;//status_reg_t'(reg2hw.status_1018.q);
  assign rcache_line[3][250].status_reg.qe    = reg2hw.status_1018.qe;
  assign rcache_line[3][250].status_reg.re    = reg2hw.status_1018.re;


  assign rcache_line[3][251].tag_reg.tag      = reg2hw.tag_1019.q;
  assign rcache_line[3][251].tag_reg.qe       = reg2hw.tag_1019.qe;
  assign rcache_line[3][251].tag_reg.re       = reg2hw.tag_1019.re;
  assign rcache_line[3][251].status_reg.status = reg2hw.status_1019.q;//status_reg_t'(reg2hw.status_1019.q);
  assign rcache_line[3][251].status_reg.qe    = reg2hw.status_1019.qe;
  assign rcache_line[3][251].status_reg.re    = reg2hw.status_1019.re;


  assign rcache_line[3][252].tag_reg.tag      = reg2hw.tag_1020.q;
  assign rcache_line[3][252].tag_reg.qe       = reg2hw.tag_1020.qe;
  assign rcache_line[3][252].tag_reg.re       = reg2hw.tag_1020.re;
  assign rcache_line[3][252].status_reg.status = reg2hw.status_1020.q;//status_reg_t'(reg2hw.status_1020.q);
  assign rcache_line[3][252].status_reg.qe    = reg2hw.status_1020.qe;
  assign rcache_line[3][252].status_reg.re    = reg2hw.status_1020.re;


  assign rcache_line[3][253].tag_reg.tag      = reg2hw.tag_1021.q;
  assign rcache_line[3][253].tag_reg.qe       = reg2hw.tag_1021.qe;
  assign rcache_line[3][253].tag_reg.re       = reg2hw.tag_1021.re;
  assign rcache_line[3][253].status_reg.status = reg2hw.status_1021.q;//status_reg_t'(reg2hw.status_1021.q);
  assign rcache_line[3][253].status_reg.qe    = reg2hw.status_1021.qe;
  assign rcache_line[3][253].status_reg.re    = reg2hw.status_1021.re;


  assign rcache_line[3][254].tag_reg.tag      = reg2hw.tag_1022.q;
  assign rcache_line[3][254].tag_reg.qe       = reg2hw.tag_1022.qe;
  assign rcache_line[3][254].tag_reg.re       = reg2hw.tag_1022.re;
  assign rcache_line[3][254].status_reg.status = reg2hw.status_1022.q;//status_reg_t'(reg2hw.status_1022.q);
  assign rcache_line[3][254].status_reg.qe    = reg2hw.status_1022.qe;
  assign rcache_line[3][254].status_reg.re    = reg2hw.status_1022.re;


  assign rcache_line[3][255].tag_reg.tag      = reg2hw.tag_1023.q;
  assign rcache_line[3][255].tag_reg.qe       = reg2hw.tag_1023.qe;
  assign rcache_line[3][255].tag_reg.re       = reg2hw.tag_1023.re;
  assign rcache_line[3][255].status_reg.status = reg2hw.status_1023.q;//status_reg_t'(reg2hw.status_1023.q);
  assign rcache_line[3][255].status_reg.qe    = reg2hw.status_1023.qe;
  assign rcache_line[3][255].status_reg.re    = reg2hw.status_1023.re;


  assign rcache_line[4][0].tag_reg.tag      = reg2hw.tag_1024.q;
  assign rcache_line[4][0].tag_reg.qe       = reg2hw.tag_1024.qe;
  assign rcache_line[4][0].tag_reg.re       = reg2hw.tag_1024.re;
  assign rcache_line[4][0].status_reg.status = reg2hw.status_1024.q;//status_reg_t'(reg2hw.status_1024.q);
  assign rcache_line[4][0].status_reg.qe    = reg2hw.status_1024.qe;
  assign rcache_line[4][0].status_reg.re    = reg2hw.status_1024.re;


  assign rcache_line[4][1].tag_reg.tag      = reg2hw.tag_1025.q;
  assign rcache_line[4][1].tag_reg.qe       = reg2hw.tag_1025.qe;
  assign rcache_line[4][1].tag_reg.re       = reg2hw.tag_1025.re;
  assign rcache_line[4][1].status_reg.status = reg2hw.status_1025.q;//status_reg_t'(reg2hw.status_1025.q);
  assign rcache_line[4][1].status_reg.qe    = reg2hw.status_1025.qe;
  assign rcache_line[4][1].status_reg.re    = reg2hw.status_1025.re;


  assign rcache_line[4][2].tag_reg.tag      = reg2hw.tag_1026.q;
  assign rcache_line[4][2].tag_reg.qe       = reg2hw.tag_1026.qe;
  assign rcache_line[4][2].tag_reg.re       = reg2hw.tag_1026.re;
  assign rcache_line[4][2].status_reg.status = reg2hw.status_1026.q;//status_reg_t'(reg2hw.status_1026.q);
  assign rcache_line[4][2].status_reg.qe    = reg2hw.status_1026.qe;
  assign rcache_line[4][2].status_reg.re    = reg2hw.status_1026.re;


  assign rcache_line[4][3].tag_reg.tag      = reg2hw.tag_1027.q;
  assign rcache_line[4][3].tag_reg.qe       = reg2hw.tag_1027.qe;
  assign rcache_line[4][3].tag_reg.re       = reg2hw.tag_1027.re;
  assign rcache_line[4][3].status_reg.status = reg2hw.status_1027.q;//status_reg_t'(reg2hw.status_1027.q);
  assign rcache_line[4][3].status_reg.qe    = reg2hw.status_1027.qe;
  assign rcache_line[4][3].status_reg.re    = reg2hw.status_1027.re;


  assign rcache_line[4][4].tag_reg.tag      = reg2hw.tag_1028.q;
  assign rcache_line[4][4].tag_reg.qe       = reg2hw.tag_1028.qe;
  assign rcache_line[4][4].tag_reg.re       = reg2hw.tag_1028.re;
  assign rcache_line[4][4].status_reg.status = reg2hw.status_1028.q;//status_reg_t'(reg2hw.status_1028.q);
  assign rcache_line[4][4].status_reg.qe    = reg2hw.status_1028.qe;
  assign rcache_line[4][4].status_reg.re    = reg2hw.status_1028.re;


  assign rcache_line[4][5].tag_reg.tag      = reg2hw.tag_1029.q;
  assign rcache_line[4][5].tag_reg.qe       = reg2hw.tag_1029.qe;
  assign rcache_line[4][5].tag_reg.re       = reg2hw.tag_1029.re;
  assign rcache_line[4][5].status_reg.status = reg2hw.status_1029.q;//status_reg_t'(reg2hw.status_1029.q);
  assign rcache_line[4][5].status_reg.qe    = reg2hw.status_1029.qe;
  assign rcache_line[4][5].status_reg.re    = reg2hw.status_1029.re;


  assign rcache_line[4][6].tag_reg.tag      = reg2hw.tag_1030.q;
  assign rcache_line[4][6].tag_reg.qe       = reg2hw.tag_1030.qe;
  assign rcache_line[4][6].tag_reg.re       = reg2hw.tag_1030.re;
  assign rcache_line[4][6].status_reg.status = reg2hw.status_1030.q;//status_reg_t'(reg2hw.status_1030.q);
  assign rcache_line[4][6].status_reg.qe    = reg2hw.status_1030.qe;
  assign rcache_line[4][6].status_reg.re    = reg2hw.status_1030.re;


  assign rcache_line[4][7].tag_reg.tag      = reg2hw.tag_1031.q;
  assign rcache_line[4][7].tag_reg.qe       = reg2hw.tag_1031.qe;
  assign rcache_line[4][7].tag_reg.re       = reg2hw.tag_1031.re;
  assign rcache_line[4][7].status_reg.status = reg2hw.status_1031.q;//status_reg_t'(reg2hw.status_1031.q);
  assign rcache_line[4][7].status_reg.qe    = reg2hw.status_1031.qe;
  assign rcache_line[4][7].status_reg.re    = reg2hw.status_1031.re;


  assign rcache_line[4][8].tag_reg.tag      = reg2hw.tag_1032.q;
  assign rcache_line[4][8].tag_reg.qe       = reg2hw.tag_1032.qe;
  assign rcache_line[4][8].tag_reg.re       = reg2hw.tag_1032.re;
  assign rcache_line[4][8].status_reg.status = reg2hw.status_1032.q;//status_reg_t'(reg2hw.status_1032.q);
  assign rcache_line[4][8].status_reg.qe    = reg2hw.status_1032.qe;
  assign rcache_line[4][8].status_reg.re    = reg2hw.status_1032.re;


  assign rcache_line[4][9].tag_reg.tag      = reg2hw.tag_1033.q;
  assign rcache_line[4][9].tag_reg.qe       = reg2hw.tag_1033.qe;
  assign rcache_line[4][9].tag_reg.re       = reg2hw.tag_1033.re;
  assign rcache_line[4][9].status_reg.status = reg2hw.status_1033.q;//status_reg_t'(reg2hw.status_1033.q);
  assign rcache_line[4][9].status_reg.qe    = reg2hw.status_1033.qe;
  assign rcache_line[4][9].status_reg.re    = reg2hw.status_1033.re;


  assign rcache_line[4][10].tag_reg.tag      = reg2hw.tag_1034.q;
  assign rcache_line[4][10].tag_reg.qe       = reg2hw.tag_1034.qe;
  assign rcache_line[4][10].tag_reg.re       = reg2hw.tag_1034.re;
  assign rcache_line[4][10].status_reg.status = reg2hw.status_1034.q;//status_reg_t'(reg2hw.status_1034.q);
  assign rcache_line[4][10].status_reg.qe    = reg2hw.status_1034.qe;
  assign rcache_line[4][10].status_reg.re    = reg2hw.status_1034.re;


  assign rcache_line[4][11].tag_reg.tag      = reg2hw.tag_1035.q;
  assign rcache_line[4][11].tag_reg.qe       = reg2hw.tag_1035.qe;
  assign rcache_line[4][11].tag_reg.re       = reg2hw.tag_1035.re;
  assign rcache_line[4][11].status_reg.status = reg2hw.status_1035.q;//status_reg_t'(reg2hw.status_1035.q);
  assign rcache_line[4][11].status_reg.qe    = reg2hw.status_1035.qe;
  assign rcache_line[4][11].status_reg.re    = reg2hw.status_1035.re;


  assign rcache_line[4][12].tag_reg.tag      = reg2hw.tag_1036.q;
  assign rcache_line[4][12].tag_reg.qe       = reg2hw.tag_1036.qe;
  assign rcache_line[4][12].tag_reg.re       = reg2hw.tag_1036.re;
  assign rcache_line[4][12].status_reg.status = reg2hw.status_1036.q;//status_reg_t'(reg2hw.status_1036.q);
  assign rcache_line[4][12].status_reg.qe    = reg2hw.status_1036.qe;
  assign rcache_line[4][12].status_reg.re    = reg2hw.status_1036.re;


  assign rcache_line[4][13].tag_reg.tag      = reg2hw.tag_1037.q;
  assign rcache_line[4][13].tag_reg.qe       = reg2hw.tag_1037.qe;
  assign rcache_line[4][13].tag_reg.re       = reg2hw.tag_1037.re;
  assign rcache_line[4][13].status_reg.status = reg2hw.status_1037.q;//status_reg_t'(reg2hw.status_1037.q);
  assign rcache_line[4][13].status_reg.qe    = reg2hw.status_1037.qe;
  assign rcache_line[4][13].status_reg.re    = reg2hw.status_1037.re;


  assign rcache_line[4][14].tag_reg.tag      = reg2hw.tag_1038.q;
  assign rcache_line[4][14].tag_reg.qe       = reg2hw.tag_1038.qe;
  assign rcache_line[4][14].tag_reg.re       = reg2hw.tag_1038.re;
  assign rcache_line[4][14].status_reg.status = reg2hw.status_1038.q;//status_reg_t'(reg2hw.status_1038.q);
  assign rcache_line[4][14].status_reg.qe    = reg2hw.status_1038.qe;
  assign rcache_line[4][14].status_reg.re    = reg2hw.status_1038.re;


  assign rcache_line[4][15].tag_reg.tag      = reg2hw.tag_1039.q;
  assign rcache_line[4][15].tag_reg.qe       = reg2hw.tag_1039.qe;
  assign rcache_line[4][15].tag_reg.re       = reg2hw.tag_1039.re;
  assign rcache_line[4][15].status_reg.status = reg2hw.status_1039.q;//status_reg_t'(reg2hw.status_1039.q);
  assign rcache_line[4][15].status_reg.qe    = reg2hw.status_1039.qe;
  assign rcache_line[4][15].status_reg.re    = reg2hw.status_1039.re;


  assign rcache_line[4][16].tag_reg.tag      = reg2hw.tag_1040.q;
  assign rcache_line[4][16].tag_reg.qe       = reg2hw.tag_1040.qe;
  assign rcache_line[4][16].tag_reg.re       = reg2hw.tag_1040.re;
  assign rcache_line[4][16].status_reg.status = reg2hw.status_1040.q;//status_reg_t'(reg2hw.status_1040.q);
  assign rcache_line[4][16].status_reg.qe    = reg2hw.status_1040.qe;
  assign rcache_line[4][16].status_reg.re    = reg2hw.status_1040.re;


  assign rcache_line[4][17].tag_reg.tag      = reg2hw.tag_1041.q;
  assign rcache_line[4][17].tag_reg.qe       = reg2hw.tag_1041.qe;
  assign rcache_line[4][17].tag_reg.re       = reg2hw.tag_1041.re;
  assign rcache_line[4][17].status_reg.status = reg2hw.status_1041.q;//status_reg_t'(reg2hw.status_1041.q);
  assign rcache_line[4][17].status_reg.qe    = reg2hw.status_1041.qe;
  assign rcache_line[4][17].status_reg.re    = reg2hw.status_1041.re;


  assign rcache_line[4][18].tag_reg.tag      = reg2hw.tag_1042.q;
  assign rcache_line[4][18].tag_reg.qe       = reg2hw.tag_1042.qe;
  assign rcache_line[4][18].tag_reg.re       = reg2hw.tag_1042.re;
  assign rcache_line[4][18].status_reg.status = reg2hw.status_1042.q;//status_reg_t'(reg2hw.status_1042.q);
  assign rcache_line[4][18].status_reg.qe    = reg2hw.status_1042.qe;
  assign rcache_line[4][18].status_reg.re    = reg2hw.status_1042.re;


  assign rcache_line[4][19].tag_reg.tag      = reg2hw.tag_1043.q;
  assign rcache_line[4][19].tag_reg.qe       = reg2hw.tag_1043.qe;
  assign rcache_line[4][19].tag_reg.re       = reg2hw.tag_1043.re;
  assign rcache_line[4][19].status_reg.status = reg2hw.status_1043.q;//status_reg_t'(reg2hw.status_1043.q);
  assign rcache_line[4][19].status_reg.qe    = reg2hw.status_1043.qe;
  assign rcache_line[4][19].status_reg.re    = reg2hw.status_1043.re;


  assign rcache_line[4][20].tag_reg.tag      = reg2hw.tag_1044.q;
  assign rcache_line[4][20].tag_reg.qe       = reg2hw.tag_1044.qe;
  assign rcache_line[4][20].tag_reg.re       = reg2hw.tag_1044.re;
  assign rcache_line[4][20].status_reg.status = reg2hw.status_1044.q;//status_reg_t'(reg2hw.status_1044.q);
  assign rcache_line[4][20].status_reg.qe    = reg2hw.status_1044.qe;
  assign rcache_line[4][20].status_reg.re    = reg2hw.status_1044.re;


  assign rcache_line[4][21].tag_reg.tag      = reg2hw.tag_1045.q;
  assign rcache_line[4][21].tag_reg.qe       = reg2hw.tag_1045.qe;
  assign rcache_line[4][21].tag_reg.re       = reg2hw.tag_1045.re;
  assign rcache_line[4][21].status_reg.status = reg2hw.status_1045.q;//status_reg_t'(reg2hw.status_1045.q);
  assign rcache_line[4][21].status_reg.qe    = reg2hw.status_1045.qe;
  assign rcache_line[4][21].status_reg.re    = reg2hw.status_1045.re;


  assign rcache_line[4][22].tag_reg.tag      = reg2hw.tag_1046.q;
  assign rcache_line[4][22].tag_reg.qe       = reg2hw.tag_1046.qe;
  assign rcache_line[4][22].tag_reg.re       = reg2hw.tag_1046.re;
  assign rcache_line[4][22].status_reg.status = reg2hw.status_1046.q;//status_reg_t'(reg2hw.status_1046.q);
  assign rcache_line[4][22].status_reg.qe    = reg2hw.status_1046.qe;
  assign rcache_line[4][22].status_reg.re    = reg2hw.status_1046.re;


  assign rcache_line[4][23].tag_reg.tag      = reg2hw.tag_1047.q;
  assign rcache_line[4][23].tag_reg.qe       = reg2hw.tag_1047.qe;
  assign rcache_line[4][23].tag_reg.re       = reg2hw.tag_1047.re;
  assign rcache_line[4][23].status_reg.status = reg2hw.status_1047.q;//status_reg_t'(reg2hw.status_1047.q);
  assign rcache_line[4][23].status_reg.qe    = reg2hw.status_1047.qe;
  assign rcache_line[4][23].status_reg.re    = reg2hw.status_1047.re;


  assign rcache_line[4][24].tag_reg.tag      = reg2hw.tag_1048.q;
  assign rcache_line[4][24].tag_reg.qe       = reg2hw.tag_1048.qe;
  assign rcache_line[4][24].tag_reg.re       = reg2hw.tag_1048.re;
  assign rcache_line[4][24].status_reg.status = reg2hw.status_1048.q;//status_reg_t'(reg2hw.status_1048.q);
  assign rcache_line[4][24].status_reg.qe    = reg2hw.status_1048.qe;
  assign rcache_line[4][24].status_reg.re    = reg2hw.status_1048.re;


  assign rcache_line[4][25].tag_reg.tag      = reg2hw.tag_1049.q;
  assign rcache_line[4][25].tag_reg.qe       = reg2hw.tag_1049.qe;
  assign rcache_line[4][25].tag_reg.re       = reg2hw.tag_1049.re;
  assign rcache_line[4][25].status_reg.status = reg2hw.status_1049.q;//status_reg_t'(reg2hw.status_1049.q);
  assign rcache_line[4][25].status_reg.qe    = reg2hw.status_1049.qe;
  assign rcache_line[4][25].status_reg.re    = reg2hw.status_1049.re;


  assign rcache_line[4][26].tag_reg.tag      = reg2hw.tag_1050.q;
  assign rcache_line[4][26].tag_reg.qe       = reg2hw.tag_1050.qe;
  assign rcache_line[4][26].tag_reg.re       = reg2hw.tag_1050.re;
  assign rcache_line[4][26].status_reg.status = reg2hw.status_1050.q;//status_reg_t'(reg2hw.status_1050.q);
  assign rcache_line[4][26].status_reg.qe    = reg2hw.status_1050.qe;
  assign rcache_line[4][26].status_reg.re    = reg2hw.status_1050.re;


  assign rcache_line[4][27].tag_reg.tag      = reg2hw.tag_1051.q;
  assign rcache_line[4][27].tag_reg.qe       = reg2hw.tag_1051.qe;
  assign rcache_line[4][27].tag_reg.re       = reg2hw.tag_1051.re;
  assign rcache_line[4][27].status_reg.status = reg2hw.status_1051.q;//status_reg_t'(reg2hw.status_1051.q);
  assign rcache_line[4][27].status_reg.qe    = reg2hw.status_1051.qe;
  assign rcache_line[4][27].status_reg.re    = reg2hw.status_1051.re;


  assign rcache_line[4][28].tag_reg.tag      = reg2hw.tag_1052.q;
  assign rcache_line[4][28].tag_reg.qe       = reg2hw.tag_1052.qe;
  assign rcache_line[4][28].tag_reg.re       = reg2hw.tag_1052.re;
  assign rcache_line[4][28].status_reg.status = reg2hw.status_1052.q;//status_reg_t'(reg2hw.status_1052.q);
  assign rcache_line[4][28].status_reg.qe    = reg2hw.status_1052.qe;
  assign rcache_line[4][28].status_reg.re    = reg2hw.status_1052.re;


  assign rcache_line[4][29].tag_reg.tag      = reg2hw.tag_1053.q;
  assign rcache_line[4][29].tag_reg.qe       = reg2hw.tag_1053.qe;
  assign rcache_line[4][29].tag_reg.re       = reg2hw.tag_1053.re;
  assign rcache_line[4][29].status_reg.status = reg2hw.status_1053.q;//status_reg_t'(reg2hw.status_1053.q);
  assign rcache_line[4][29].status_reg.qe    = reg2hw.status_1053.qe;
  assign rcache_line[4][29].status_reg.re    = reg2hw.status_1053.re;


  assign rcache_line[4][30].tag_reg.tag      = reg2hw.tag_1054.q;
  assign rcache_line[4][30].tag_reg.qe       = reg2hw.tag_1054.qe;
  assign rcache_line[4][30].tag_reg.re       = reg2hw.tag_1054.re;
  assign rcache_line[4][30].status_reg.status = reg2hw.status_1054.q;//status_reg_t'(reg2hw.status_1054.q);
  assign rcache_line[4][30].status_reg.qe    = reg2hw.status_1054.qe;
  assign rcache_line[4][30].status_reg.re    = reg2hw.status_1054.re;


  assign rcache_line[4][31].tag_reg.tag      = reg2hw.tag_1055.q;
  assign rcache_line[4][31].tag_reg.qe       = reg2hw.tag_1055.qe;
  assign rcache_line[4][31].tag_reg.re       = reg2hw.tag_1055.re;
  assign rcache_line[4][31].status_reg.status = reg2hw.status_1055.q;//status_reg_t'(reg2hw.status_1055.q);
  assign rcache_line[4][31].status_reg.qe    = reg2hw.status_1055.qe;
  assign rcache_line[4][31].status_reg.re    = reg2hw.status_1055.re;


  assign rcache_line[4][32].tag_reg.tag      = reg2hw.tag_1056.q;
  assign rcache_line[4][32].tag_reg.qe       = reg2hw.tag_1056.qe;
  assign rcache_line[4][32].tag_reg.re       = reg2hw.tag_1056.re;
  assign rcache_line[4][32].status_reg.status = reg2hw.status_1056.q;//status_reg_t'(reg2hw.status_1056.q);
  assign rcache_line[4][32].status_reg.qe    = reg2hw.status_1056.qe;
  assign rcache_line[4][32].status_reg.re    = reg2hw.status_1056.re;


  assign rcache_line[4][33].tag_reg.tag      = reg2hw.tag_1057.q;
  assign rcache_line[4][33].tag_reg.qe       = reg2hw.tag_1057.qe;
  assign rcache_line[4][33].tag_reg.re       = reg2hw.tag_1057.re;
  assign rcache_line[4][33].status_reg.status = reg2hw.status_1057.q;//status_reg_t'(reg2hw.status_1057.q);
  assign rcache_line[4][33].status_reg.qe    = reg2hw.status_1057.qe;
  assign rcache_line[4][33].status_reg.re    = reg2hw.status_1057.re;


  assign rcache_line[4][34].tag_reg.tag      = reg2hw.tag_1058.q;
  assign rcache_line[4][34].tag_reg.qe       = reg2hw.tag_1058.qe;
  assign rcache_line[4][34].tag_reg.re       = reg2hw.tag_1058.re;
  assign rcache_line[4][34].status_reg.status = reg2hw.status_1058.q;//status_reg_t'(reg2hw.status_1058.q);
  assign rcache_line[4][34].status_reg.qe    = reg2hw.status_1058.qe;
  assign rcache_line[4][34].status_reg.re    = reg2hw.status_1058.re;


  assign rcache_line[4][35].tag_reg.tag      = reg2hw.tag_1059.q;
  assign rcache_line[4][35].tag_reg.qe       = reg2hw.tag_1059.qe;
  assign rcache_line[4][35].tag_reg.re       = reg2hw.tag_1059.re;
  assign rcache_line[4][35].status_reg.status = reg2hw.status_1059.q;//status_reg_t'(reg2hw.status_1059.q);
  assign rcache_line[4][35].status_reg.qe    = reg2hw.status_1059.qe;
  assign rcache_line[4][35].status_reg.re    = reg2hw.status_1059.re;


  assign rcache_line[4][36].tag_reg.tag      = reg2hw.tag_1060.q;
  assign rcache_line[4][36].tag_reg.qe       = reg2hw.tag_1060.qe;
  assign rcache_line[4][36].tag_reg.re       = reg2hw.tag_1060.re;
  assign rcache_line[4][36].status_reg.status = reg2hw.status_1060.q;//status_reg_t'(reg2hw.status_1060.q);
  assign rcache_line[4][36].status_reg.qe    = reg2hw.status_1060.qe;
  assign rcache_line[4][36].status_reg.re    = reg2hw.status_1060.re;


  assign rcache_line[4][37].tag_reg.tag      = reg2hw.tag_1061.q;
  assign rcache_line[4][37].tag_reg.qe       = reg2hw.tag_1061.qe;
  assign rcache_line[4][37].tag_reg.re       = reg2hw.tag_1061.re;
  assign rcache_line[4][37].status_reg.status = reg2hw.status_1061.q;//status_reg_t'(reg2hw.status_1061.q);
  assign rcache_line[4][37].status_reg.qe    = reg2hw.status_1061.qe;
  assign rcache_line[4][37].status_reg.re    = reg2hw.status_1061.re;


  assign rcache_line[4][38].tag_reg.tag      = reg2hw.tag_1062.q;
  assign rcache_line[4][38].tag_reg.qe       = reg2hw.tag_1062.qe;
  assign rcache_line[4][38].tag_reg.re       = reg2hw.tag_1062.re;
  assign rcache_line[4][38].status_reg.status = reg2hw.status_1062.q;//status_reg_t'(reg2hw.status_1062.q);
  assign rcache_line[4][38].status_reg.qe    = reg2hw.status_1062.qe;
  assign rcache_line[4][38].status_reg.re    = reg2hw.status_1062.re;


  assign rcache_line[4][39].tag_reg.tag      = reg2hw.tag_1063.q;
  assign rcache_line[4][39].tag_reg.qe       = reg2hw.tag_1063.qe;
  assign rcache_line[4][39].tag_reg.re       = reg2hw.tag_1063.re;
  assign rcache_line[4][39].status_reg.status = reg2hw.status_1063.q;//status_reg_t'(reg2hw.status_1063.q);
  assign rcache_line[4][39].status_reg.qe    = reg2hw.status_1063.qe;
  assign rcache_line[4][39].status_reg.re    = reg2hw.status_1063.re;


  assign rcache_line[4][40].tag_reg.tag      = reg2hw.tag_1064.q;
  assign rcache_line[4][40].tag_reg.qe       = reg2hw.tag_1064.qe;
  assign rcache_line[4][40].tag_reg.re       = reg2hw.tag_1064.re;
  assign rcache_line[4][40].status_reg.status = reg2hw.status_1064.q;//status_reg_t'(reg2hw.status_1064.q);
  assign rcache_line[4][40].status_reg.qe    = reg2hw.status_1064.qe;
  assign rcache_line[4][40].status_reg.re    = reg2hw.status_1064.re;


  assign rcache_line[4][41].tag_reg.tag      = reg2hw.tag_1065.q;
  assign rcache_line[4][41].tag_reg.qe       = reg2hw.tag_1065.qe;
  assign rcache_line[4][41].tag_reg.re       = reg2hw.tag_1065.re;
  assign rcache_line[4][41].status_reg.status = reg2hw.status_1065.q;//status_reg_t'(reg2hw.status_1065.q);
  assign rcache_line[4][41].status_reg.qe    = reg2hw.status_1065.qe;
  assign rcache_line[4][41].status_reg.re    = reg2hw.status_1065.re;


  assign rcache_line[4][42].tag_reg.tag      = reg2hw.tag_1066.q;
  assign rcache_line[4][42].tag_reg.qe       = reg2hw.tag_1066.qe;
  assign rcache_line[4][42].tag_reg.re       = reg2hw.tag_1066.re;
  assign rcache_line[4][42].status_reg.status = reg2hw.status_1066.q;//status_reg_t'(reg2hw.status_1066.q);
  assign rcache_line[4][42].status_reg.qe    = reg2hw.status_1066.qe;
  assign rcache_line[4][42].status_reg.re    = reg2hw.status_1066.re;


  assign rcache_line[4][43].tag_reg.tag      = reg2hw.tag_1067.q;
  assign rcache_line[4][43].tag_reg.qe       = reg2hw.tag_1067.qe;
  assign rcache_line[4][43].tag_reg.re       = reg2hw.tag_1067.re;
  assign rcache_line[4][43].status_reg.status = reg2hw.status_1067.q;//status_reg_t'(reg2hw.status_1067.q);
  assign rcache_line[4][43].status_reg.qe    = reg2hw.status_1067.qe;
  assign rcache_line[4][43].status_reg.re    = reg2hw.status_1067.re;


  assign rcache_line[4][44].tag_reg.tag      = reg2hw.tag_1068.q;
  assign rcache_line[4][44].tag_reg.qe       = reg2hw.tag_1068.qe;
  assign rcache_line[4][44].tag_reg.re       = reg2hw.tag_1068.re;
  assign rcache_line[4][44].status_reg.status = reg2hw.status_1068.q;//status_reg_t'(reg2hw.status_1068.q);
  assign rcache_line[4][44].status_reg.qe    = reg2hw.status_1068.qe;
  assign rcache_line[4][44].status_reg.re    = reg2hw.status_1068.re;


  assign rcache_line[4][45].tag_reg.tag      = reg2hw.tag_1069.q;
  assign rcache_line[4][45].tag_reg.qe       = reg2hw.tag_1069.qe;
  assign rcache_line[4][45].tag_reg.re       = reg2hw.tag_1069.re;
  assign rcache_line[4][45].status_reg.status = reg2hw.status_1069.q;//status_reg_t'(reg2hw.status_1069.q);
  assign rcache_line[4][45].status_reg.qe    = reg2hw.status_1069.qe;
  assign rcache_line[4][45].status_reg.re    = reg2hw.status_1069.re;


  assign rcache_line[4][46].tag_reg.tag      = reg2hw.tag_1070.q;
  assign rcache_line[4][46].tag_reg.qe       = reg2hw.tag_1070.qe;
  assign rcache_line[4][46].tag_reg.re       = reg2hw.tag_1070.re;
  assign rcache_line[4][46].status_reg.status = reg2hw.status_1070.q;//status_reg_t'(reg2hw.status_1070.q);
  assign rcache_line[4][46].status_reg.qe    = reg2hw.status_1070.qe;
  assign rcache_line[4][46].status_reg.re    = reg2hw.status_1070.re;


  assign rcache_line[4][47].tag_reg.tag      = reg2hw.tag_1071.q;
  assign rcache_line[4][47].tag_reg.qe       = reg2hw.tag_1071.qe;
  assign rcache_line[4][47].tag_reg.re       = reg2hw.tag_1071.re;
  assign rcache_line[4][47].status_reg.status = reg2hw.status_1071.q;//status_reg_t'(reg2hw.status_1071.q);
  assign rcache_line[4][47].status_reg.qe    = reg2hw.status_1071.qe;
  assign rcache_line[4][47].status_reg.re    = reg2hw.status_1071.re;


  assign rcache_line[4][48].tag_reg.tag      = reg2hw.tag_1072.q;
  assign rcache_line[4][48].tag_reg.qe       = reg2hw.tag_1072.qe;
  assign rcache_line[4][48].tag_reg.re       = reg2hw.tag_1072.re;
  assign rcache_line[4][48].status_reg.status = reg2hw.status_1072.q;//status_reg_t'(reg2hw.status_1072.q);
  assign rcache_line[4][48].status_reg.qe    = reg2hw.status_1072.qe;
  assign rcache_line[4][48].status_reg.re    = reg2hw.status_1072.re;


  assign rcache_line[4][49].tag_reg.tag      = reg2hw.tag_1073.q;
  assign rcache_line[4][49].tag_reg.qe       = reg2hw.tag_1073.qe;
  assign rcache_line[4][49].tag_reg.re       = reg2hw.tag_1073.re;
  assign rcache_line[4][49].status_reg.status = reg2hw.status_1073.q;//status_reg_t'(reg2hw.status_1073.q);
  assign rcache_line[4][49].status_reg.qe    = reg2hw.status_1073.qe;
  assign rcache_line[4][49].status_reg.re    = reg2hw.status_1073.re;


  assign rcache_line[4][50].tag_reg.tag      = reg2hw.tag_1074.q;
  assign rcache_line[4][50].tag_reg.qe       = reg2hw.tag_1074.qe;
  assign rcache_line[4][50].tag_reg.re       = reg2hw.tag_1074.re;
  assign rcache_line[4][50].status_reg.status = reg2hw.status_1074.q;//status_reg_t'(reg2hw.status_1074.q);
  assign rcache_line[4][50].status_reg.qe    = reg2hw.status_1074.qe;
  assign rcache_line[4][50].status_reg.re    = reg2hw.status_1074.re;


  assign rcache_line[4][51].tag_reg.tag      = reg2hw.tag_1075.q;
  assign rcache_line[4][51].tag_reg.qe       = reg2hw.tag_1075.qe;
  assign rcache_line[4][51].tag_reg.re       = reg2hw.tag_1075.re;
  assign rcache_line[4][51].status_reg.status = reg2hw.status_1075.q;//status_reg_t'(reg2hw.status_1075.q);
  assign rcache_line[4][51].status_reg.qe    = reg2hw.status_1075.qe;
  assign rcache_line[4][51].status_reg.re    = reg2hw.status_1075.re;


  assign rcache_line[4][52].tag_reg.tag      = reg2hw.tag_1076.q;
  assign rcache_line[4][52].tag_reg.qe       = reg2hw.tag_1076.qe;
  assign rcache_line[4][52].tag_reg.re       = reg2hw.tag_1076.re;
  assign rcache_line[4][52].status_reg.status = reg2hw.status_1076.q;//status_reg_t'(reg2hw.status_1076.q);
  assign rcache_line[4][52].status_reg.qe    = reg2hw.status_1076.qe;
  assign rcache_line[4][52].status_reg.re    = reg2hw.status_1076.re;


  assign rcache_line[4][53].tag_reg.tag      = reg2hw.tag_1077.q;
  assign rcache_line[4][53].tag_reg.qe       = reg2hw.tag_1077.qe;
  assign rcache_line[4][53].tag_reg.re       = reg2hw.tag_1077.re;
  assign rcache_line[4][53].status_reg.status = reg2hw.status_1077.q;//status_reg_t'(reg2hw.status_1077.q);
  assign rcache_line[4][53].status_reg.qe    = reg2hw.status_1077.qe;
  assign rcache_line[4][53].status_reg.re    = reg2hw.status_1077.re;


  assign rcache_line[4][54].tag_reg.tag      = reg2hw.tag_1078.q;
  assign rcache_line[4][54].tag_reg.qe       = reg2hw.tag_1078.qe;
  assign rcache_line[4][54].tag_reg.re       = reg2hw.tag_1078.re;
  assign rcache_line[4][54].status_reg.status = reg2hw.status_1078.q;//status_reg_t'(reg2hw.status_1078.q);
  assign rcache_line[4][54].status_reg.qe    = reg2hw.status_1078.qe;
  assign rcache_line[4][54].status_reg.re    = reg2hw.status_1078.re;


  assign rcache_line[4][55].tag_reg.tag      = reg2hw.tag_1079.q;
  assign rcache_line[4][55].tag_reg.qe       = reg2hw.tag_1079.qe;
  assign rcache_line[4][55].tag_reg.re       = reg2hw.tag_1079.re;
  assign rcache_line[4][55].status_reg.status = reg2hw.status_1079.q;//status_reg_t'(reg2hw.status_1079.q);
  assign rcache_line[4][55].status_reg.qe    = reg2hw.status_1079.qe;
  assign rcache_line[4][55].status_reg.re    = reg2hw.status_1079.re;


  assign rcache_line[4][56].tag_reg.tag      = reg2hw.tag_1080.q;
  assign rcache_line[4][56].tag_reg.qe       = reg2hw.tag_1080.qe;
  assign rcache_line[4][56].tag_reg.re       = reg2hw.tag_1080.re;
  assign rcache_line[4][56].status_reg.status = reg2hw.status_1080.q;//status_reg_t'(reg2hw.status_1080.q);
  assign rcache_line[4][56].status_reg.qe    = reg2hw.status_1080.qe;
  assign rcache_line[4][56].status_reg.re    = reg2hw.status_1080.re;


  assign rcache_line[4][57].tag_reg.tag      = reg2hw.tag_1081.q;
  assign rcache_line[4][57].tag_reg.qe       = reg2hw.tag_1081.qe;
  assign rcache_line[4][57].tag_reg.re       = reg2hw.tag_1081.re;
  assign rcache_line[4][57].status_reg.status = reg2hw.status_1081.q;//status_reg_t'(reg2hw.status_1081.q);
  assign rcache_line[4][57].status_reg.qe    = reg2hw.status_1081.qe;
  assign rcache_line[4][57].status_reg.re    = reg2hw.status_1081.re;


  assign rcache_line[4][58].tag_reg.tag      = reg2hw.tag_1082.q;
  assign rcache_line[4][58].tag_reg.qe       = reg2hw.tag_1082.qe;
  assign rcache_line[4][58].tag_reg.re       = reg2hw.tag_1082.re;
  assign rcache_line[4][58].status_reg.status = reg2hw.status_1082.q;//status_reg_t'(reg2hw.status_1082.q);
  assign rcache_line[4][58].status_reg.qe    = reg2hw.status_1082.qe;
  assign rcache_line[4][58].status_reg.re    = reg2hw.status_1082.re;


  assign rcache_line[4][59].tag_reg.tag      = reg2hw.tag_1083.q;
  assign rcache_line[4][59].tag_reg.qe       = reg2hw.tag_1083.qe;
  assign rcache_line[4][59].tag_reg.re       = reg2hw.tag_1083.re;
  assign rcache_line[4][59].status_reg.status = reg2hw.status_1083.q;//status_reg_t'(reg2hw.status_1083.q);
  assign rcache_line[4][59].status_reg.qe    = reg2hw.status_1083.qe;
  assign rcache_line[4][59].status_reg.re    = reg2hw.status_1083.re;


  assign rcache_line[4][60].tag_reg.tag      = reg2hw.tag_1084.q;
  assign rcache_line[4][60].tag_reg.qe       = reg2hw.tag_1084.qe;
  assign rcache_line[4][60].tag_reg.re       = reg2hw.tag_1084.re;
  assign rcache_line[4][60].status_reg.status = reg2hw.status_1084.q;//status_reg_t'(reg2hw.status_1084.q);
  assign rcache_line[4][60].status_reg.qe    = reg2hw.status_1084.qe;
  assign rcache_line[4][60].status_reg.re    = reg2hw.status_1084.re;


  assign rcache_line[4][61].tag_reg.tag      = reg2hw.tag_1085.q;
  assign rcache_line[4][61].tag_reg.qe       = reg2hw.tag_1085.qe;
  assign rcache_line[4][61].tag_reg.re       = reg2hw.tag_1085.re;
  assign rcache_line[4][61].status_reg.status = reg2hw.status_1085.q;//status_reg_t'(reg2hw.status_1085.q);
  assign rcache_line[4][61].status_reg.qe    = reg2hw.status_1085.qe;
  assign rcache_line[4][61].status_reg.re    = reg2hw.status_1085.re;


  assign rcache_line[4][62].tag_reg.tag      = reg2hw.tag_1086.q;
  assign rcache_line[4][62].tag_reg.qe       = reg2hw.tag_1086.qe;
  assign rcache_line[4][62].tag_reg.re       = reg2hw.tag_1086.re;
  assign rcache_line[4][62].status_reg.status = reg2hw.status_1086.q;//status_reg_t'(reg2hw.status_1086.q);
  assign rcache_line[4][62].status_reg.qe    = reg2hw.status_1086.qe;
  assign rcache_line[4][62].status_reg.re    = reg2hw.status_1086.re;


  assign rcache_line[4][63].tag_reg.tag      = reg2hw.tag_1087.q;
  assign rcache_line[4][63].tag_reg.qe       = reg2hw.tag_1087.qe;
  assign rcache_line[4][63].tag_reg.re       = reg2hw.tag_1087.re;
  assign rcache_line[4][63].status_reg.status = reg2hw.status_1087.q;//status_reg_t'(reg2hw.status_1087.q);
  assign rcache_line[4][63].status_reg.qe    = reg2hw.status_1087.qe;
  assign rcache_line[4][63].status_reg.re    = reg2hw.status_1087.re;


  assign rcache_line[4][64].tag_reg.tag      = reg2hw.tag_1088.q;
  assign rcache_line[4][64].tag_reg.qe       = reg2hw.tag_1088.qe;
  assign rcache_line[4][64].tag_reg.re       = reg2hw.tag_1088.re;
  assign rcache_line[4][64].status_reg.status = reg2hw.status_1088.q;//status_reg_t'(reg2hw.status_1088.q);
  assign rcache_line[4][64].status_reg.qe    = reg2hw.status_1088.qe;
  assign rcache_line[4][64].status_reg.re    = reg2hw.status_1088.re;


  assign rcache_line[4][65].tag_reg.tag      = reg2hw.tag_1089.q;
  assign rcache_line[4][65].tag_reg.qe       = reg2hw.tag_1089.qe;
  assign rcache_line[4][65].tag_reg.re       = reg2hw.tag_1089.re;
  assign rcache_line[4][65].status_reg.status = reg2hw.status_1089.q;//status_reg_t'(reg2hw.status_1089.q);
  assign rcache_line[4][65].status_reg.qe    = reg2hw.status_1089.qe;
  assign rcache_line[4][65].status_reg.re    = reg2hw.status_1089.re;


  assign rcache_line[4][66].tag_reg.tag      = reg2hw.tag_1090.q;
  assign rcache_line[4][66].tag_reg.qe       = reg2hw.tag_1090.qe;
  assign rcache_line[4][66].tag_reg.re       = reg2hw.tag_1090.re;
  assign rcache_line[4][66].status_reg.status = reg2hw.status_1090.q;//status_reg_t'(reg2hw.status_1090.q);
  assign rcache_line[4][66].status_reg.qe    = reg2hw.status_1090.qe;
  assign rcache_line[4][66].status_reg.re    = reg2hw.status_1090.re;


  assign rcache_line[4][67].tag_reg.tag      = reg2hw.tag_1091.q;
  assign rcache_line[4][67].tag_reg.qe       = reg2hw.tag_1091.qe;
  assign rcache_line[4][67].tag_reg.re       = reg2hw.tag_1091.re;
  assign rcache_line[4][67].status_reg.status = reg2hw.status_1091.q;//status_reg_t'(reg2hw.status_1091.q);
  assign rcache_line[4][67].status_reg.qe    = reg2hw.status_1091.qe;
  assign rcache_line[4][67].status_reg.re    = reg2hw.status_1091.re;


  assign rcache_line[4][68].tag_reg.tag      = reg2hw.tag_1092.q;
  assign rcache_line[4][68].tag_reg.qe       = reg2hw.tag_1092.qe;
  assign rcache_line[4][68].tag_reg.re       = reg2hw.tag_1092.re;
  assign rcache_line[4][68].status_reg.status = reg2hw.status_1092.q;//status_reg_t'(reg2hw.status_1092.q);
  assign rcache_line[4][68].status_reg.qe    = reg2hw.status_1092.qe;
  assign rcache_line[4][68].status_reg.re    = reg2hw.status_1092.re;


  assign rcache_line[4][69].tag_reg.tag      = reg2hw.tag_1093.q;
  assign rcache_line[4][69].tag_reg.qe       = reg2hw.tag_1093.qe;
  assign rcache_line[4][69].tag_reg.re       = reg2hw.tag_1093.re;
  assign rcache_line[4][69].status_reg.status = reg2hw.status_1093.q;//status_reg_t'(reg2hw.status_1093.q);
  assign rcache_line[4][69].status_reg.qe    = reg2hw.status_1093.qe;
  assign rcache_line[4][69].status_reg.re    = reg2hw.status_1093.re;


  assign rcache_line[4][70].tag_reg.tag      = reg2hw.tag_1094.q;
  assign rcache_line[4][70].tag_reg.qe       = reg2hw.tag_1094.qe;
  assign rcache_line[4][70].tag_reg.re       = reg2hw.tag_1094.re;
  assign rcache_line[4][70].status_reg.status = reg2hw.status_1094.q;//status_reg_t'(reg2hw.status_1094.q);
  assign rcache_line[4][70].status_reg.qe    = reg2hw.status_1094.qe;
  assign rcache_line[4][70].status_reg.re    = reg2hw.status_1094.re;


  assign rcache_line[4][71].tag_reg.tag      = reg2hw.tag_1095.q;
  assign rcache_line[4][71].tag_reg.qe       = reg2hw.tag_1095.qe;
  assign rcache_line[4][71].tag_reg.re       = reg2hw.tag_1095.re;
  assign rcache_line[4][71].status_reg.status = reg2hw.status_1095.q;//status_reg_t'(reg2hw.status_1095.q);
  assign rcache_line[4][71].status_reg.qe    = reg2hw.status_1095.qe;
  assign rcache_line[4][71].status_reg.re    = reg2hw.status_1095.re;


  assign rcache_line[4][72].tag_reg.tag      = reg2hw.tag_1096.q;
  assign rcache_line[4][72].tag_reg.qe       = reg2hw.tag_1096.qe;
  assign rcache_line[4][72].tag_reg.re       = reg2hw.tag_1096.re;
  assign rcache_line[4][72].status_reg.status = reg2hw.status_1096.q;//status_reg_t'(reg2hw.status_1096.q);
  assign rcache_line[4][72].status_reg.qe    = reg2hw.status_1096.qe;
  assign rcache_line[4][72].status_reg.re    = reg2hw.status_1096.re;


  assign rcache_line[4][73].tag_reg.tag      = reg2hw.tag_1097.q;
  assign rcache_line[4][73].tag_reg.qe       = reg2hw.tag_1097.qe;
  assign rcache_line[4][73].tag_reg.re       = reg2hw.tag_1097.re;
  assign rcache_line[4][73].status_reg.status = reg2hw.status_1097.q;//status_reg_t'(reg2hw.status_1097.q);
  assign rcache_line[4][73].status_reg.qe    = reg2hw.status_1097.qe;
  assign rcache_line[4][73].status_reg.re    = reg2hw.status_1097.re;


  assign rcache_line[4][74].tag_reg.tag      = reg2hw.tag_1098.q;
  assign rcache_line[4][74].tag_reg.qe       = reg2hw.tag_1098.qe;
  assign rcache_line[4][74].tag_reg.re       = reg2hw.tag_1098.re;
  assign rcache_line[4][74].status_reg.status = reg2hw.status_1098.q;//status_reg_t'(reg2hw.status_1098.q);
  assign rcache_line[4][74].status_reg.qe    = reg2hw.status_1098.qe;
  assign rcache_line[4][74].status_reg.re    = reg2hw.status_1098.re;


  assign rcache_line[4][75].tag_reg.tag      = reg2hw.tag_1099.q;
  assign rcache_line[4][75].tag_reg.qe       = reg2hw.tag_1099.qe;
  assign rcache_line[4][75].tag_reg.re       = reg2hw.tag_1099.re;
  assign rcache_line[4][75].status_reg.status = reg2hw.status_1099.q;//status_reg_t'(reg2hw.status_1099.q);
  assign rcache_line[4][75].status_reg.qe    = reg2hw.status_1099.qe;
  assign rcache_line[4][75].status_reg.re    = reg2hw.status_1099.re;


  assign rcache_line[4][76].tag_reg.tag      = reg2hw.tag_1100.q;
  assign rcache_line[4][76].tag_reg.qe       = reg2hw.tag_1100.qe;
  assign rcache_line[4][76].tag_reg.re       = reg2hw.tag_1100.re;
  assign rcache_line[4][76].status_reg.status = reg2hw.status_1100.q;//status_reg_t'(reg2hw.status_1100.q);
  assign rcache_line[4][76].status_reg.qe    = reg2hw.status_1100.qe;
  assign rcache_line[4][76].status_reg.re    = reg2hw.status_1100.re;


  assign rcache_line[4][77].tag_reg.tag      = reg2hw.tag_1101.q;
  assign rcache_line[4][77].tag_reg.qe       = reg2hw.tag_1101.qe;
  assign rcache_line[4][77].tag_reg.re       = reg2hw.tag_1101.re;
  assign rcache_line[4][77].status_reg.status = reg2hw.status_1101.q;//status_reg_t'(reg2hw.status_1101.q);
  assign rcache_line[4][77].status_reg.qe    = reg2hw.status_1101.qe;
  assign rcache_line[4][77].status_reg.re    = reg2hw.status_1101.re;


  assign rcache_line[4][78].tag_reg.tag      = reg2hw.tag_1102.q;
  assign rcache_line[4][78].tag_reg.qe       = reg2hw.tag_1102.qe;
  assign rcache_line[4][78].tag_reg.re       = reg2hw.tag_1102.re;
  assign rcache_line[4][78].status_reg.status = reg2hw.status_1102.q;//status_reg_t'(reg2hw.status_1102.q);
  assign rcache_line[4][78].status_reg.qe    = reg2hw.status_1102.qe;
  assign rcache_line[4][78].status_reg.re    = reg2hw.status_1102.re;


  assign rcache_line[4][79].tag_reg.tag      = reg2hw.tag_1103.q;
  assign rcache_line[4][79].tag_reg.qe       = reg2hw.tag_1103.qe;
  assign rcache_line[4][79].tag_reg.re       = reg2hw.tag_1103.re;
  assign rcache_line[4][79].status_reg.status = reg2hw.status_1103.q;//status_reg_t'(reg2hw.status_1103.q);
  assign rcache_line[4][79].status_reg.qe    = reg2hw.status_1103.qe;
  assign rcache_line[4][79].status_reg.re    = reg2hw.status_1103.re;


  assign rcache_line[4][80].tag_reg.tag      = reg2hw.tag_1104.q;
  assign rcache_line[4][80].tag_reg.qe       = reg2hw.tag_1104.qe;
  assign rcache_line[4][80].tag_reg.re       = reg2hw.tag_1104.re;
  assign rcache_line[4][80].status_reg.status = reg2hw.status_1104.q;//status_reg_t'(reg2hw.status_1104.q);
  assign rcache_line[4][80].status_reg.qe    = reg2hw.status_1104.qe;
  assign rcache_line[4][80].status_reg.re    = reg2hw.status_1104.re;


  assign rcache_line[4][81].tag_reg.tag      = reg2hw.tag_1105.q;
  assign rcache_line[4][81].tag_reg.qe       = reg2hw.tag_1105.qe;
  assign rcache_line[4][81].tag_reg.re       = reg2hw.tag_1105.re;
  assign rcache_line[4][81].status_reg.status = reg2hw.status_1105.q;//status_reg_t'(reg2hw.status_1105.q);
  assign rcache_line[4][81].status_reg.qe    = reg2hw.status_1105.qe;
  assign rcache_line[4][81].status_reg.re    = reg2hw.status_1105.re;


  assign rcache_line[4][82].tag_reg.tag      = reg2hw.tag_1106.q;
  assign rcache_line[4][82].tag_reg.qe       = reg2hw.tag_1106.qe;
  assign rcache_line[4][82].tag_reg.re       = reg2hw.tag_1106.re;
  assign rcache_line[4][82].status_reg.status = reg2hw.status_1106.q;//status_reg_t'(reg2hw.status_1106.q);
  assign rcache_line[4][82].status_reg.qe    = reg2hw.status_1106.qe;
  assign rcache_line[4][82].status_reg.re    = reg2hw.status_1106.re;


  assign rcache_line[4][83].tag_reg.tag      = reg2hw.tag_1107.q;
  assign rcache_line[4][83].tag_reg.qe       = reg2hw.tag_1107.qe;
  assign rcache_line[4][83].tag_reg.re       = reg2hw.tag_1107.re;
  assign rcache_line[4][83].status_reg.status = reg2hw.status_1107.q;//status_reg_t'(reg2hw.status_1107.q);
  assign rcache_line[4][83].status_reg.qe    = reg2hw.status_1107.qe;
  assign rcache_line[4][83].status_reg.re    = reg2hw.status_1107.re;


  assign rcache_line[4][84].tag_reg.tag      = reg2hw.tag_1108.q;
  assign rcache_line[4][84].tag_reg.qe       = reg2hw.tag_1108.qe;
  assign rcache_line[4][84].tag_reg.re       = reg2hw.tag_1108.re;
  assign rcache_line[4][84].status_reg.status = reg2hw.status_1108.q;//status_reg_t'(reg2hw.status_1108.q);
  assign rcache_line[4][84].status_reg.qe    = reg2hw.status_1108.qe;
  assign rcache_line[4][84].status_reg.re    = reg2hw.status_1108.re;


  assign rcache_line[4][85].tag_reg.tag      = reg2hw.tag_1109.q;
  assign rcache_line[4][85].tag_reg.qe       = reg2hw.tag_1109.qe;
  assign rcache_line[4][85].tag_reg.re       = reg2hw.tag_1109.re;
  assign rcache_line[4][85].status_reg.status = reg2hw.status_1109.q;//status_reg_t'(reg2hw.status_1109.q);
  assign rcache_line[4][85].status_reg.qe    = reg2hw.status_1109.qe;
  assign rcache_line[4][85].status_reg.re    = reg2hw.status_1109.re;


  assign rcache_line[4][86].tag_reg.tag      = reg2hw.tag_1110.q;
  assign rcache_line[4][86].tag_reg.qe       = reg2hw.tag_1110.qe;
  assign rcache_line[4][86].tag_reg.re       = reg2hw.tag_1110.re;
  assign rcache_line[4][86].status_reg.status = reg2hw.status_1110.q;//status_reg_t'(reg2hw.status_1110.q);
  assign rcache_line[4][86].status_reg.qe    = reg2hw.status_1110.qe;
  assign rcache_line[4][86].status_reg.re    = reg2hw.status_1110.re;


  assign rcache_line[4][87].tag_reg.tag      = reg2hw.tag_1111.q;
  assign rcache_line[4][87].tag_reg.qe       = reg2hw.tag_1111.qe;
  assign rcache_line[4][87].tag_reg.re       = reg2hw.tag_1111.re;
  assign rcache_line[4][87].status_reg.status = reg2hw.status_1111.q;//status_reg_t'(reg2hw.status_1111.q);
  assign rcache_line[4][87].status_reg.qe    = reg2hw.status_1111.qe;
  assign rcache_line[4][87].status_reg.re    = reg2hw.status_1111.re;


  assign rcache_line[4][88].tag_reg.tag      = reg2hw.tag_1112.q;
  assign rcache_line[4][88].tag_reg.qe       = reg2hw.tag_1112.qe;
  assign rcache_line[4][88].tag_reg.re       = reg2hw.tag_1112.re;
  assign rcache_line[4][88].status_reg.status = reg2hw.status_1112.q;//status_reg_t'(reg2hw.status_1112.q);
  assign rcache_line[4][88].status_reg.qe    = reg2hw.status_1112.qe;
  assign rcache_line[4][88].status_reg.re    = reg2hw.status_1112.re;


  assign rcache_line[4][89].tag_reg.tag      = reg2hw.tag_1113.q;
  assign rcache_line[4][89].tag_reg.qe       = reg2hw.tag_1113.qe;
  assign rcache_line[4][89].tag_reg.re       = reg2hw.tag_1113.re;
  assign rcache_line[4][89].status_reg.status = reg2hw.status_1113.q;//status_reg_t'(reg2hw.status_1113.q);
  assign rcache_line[4][89].status_reg.qe    = reg2hw.status_1113.qe;
  assign rcache_line[4][89].status_reg.re    = reg2hw.status_1113.re;


  assign rcache_line[4][90].tag_reg.tag      = reg2hw.tag_1114.q;
  assign rcache_line[4][90].tag_reg.qe       = reg2hw.tag_1114.qe;
  assign rcache_line[4][90].tag_reg.re       = reg2hw.tag_1114.re;
  assign rcache_line[4][90].status_reg.status = reg2hw.status_1114.q;//status_reg_t'(reg2hw.status_1114.q);
  assign rcache_line[4][90].status_reg.qe    = reg2hw.status_1114.qe;
  assign rcache_line[4][90].status_reg.re    = reg2hw.status_1114.re;


  assign rcache_line[4][91].tag_reg.tag      = reg2hw.tag_1115.q;
  assign rcache_line[4][91].tag_reg.qe       = reg2hw.tag_1115.qe;
  assign rcache_line[4][91].tag_reg.re       = reg2hw.tag_1115.re;
  assign rcache_line[4][91].status_reg.status = reg2hw.status_1115.q;//status_reg_t'(reg2hw.status_1115.q);
  assign rcache_line[4][91].status_reg.qe    = reg2hw.status_1115.qe;
  assign rcache_line[4][91].status_reg.re    = reg2hw.status_1115.re;


  assign rcache_line[4][92].tag_reg.tag      = reg2hw.tag_1116.q;
  assign rcache_line[4][92].tag_reg.qe       = reg2hw.tag_1116.qe;
  assign rcache_line[4][92].tag_reg.re       = reg2hw.tag_1116.re;
  assign rcache_line[4][92].status_reg.status = reg2hw.status_1116.q;//status_reg_t'(reg2hw.status_1116.q);
  assign rcache_line[4][92].status_reg.qe    = reg2hw.status_1116.qe;
  assign rcache_line[4][92].status_reg.re    = reg2hw.status_1116.re;


  assign rcache_line[4][93].tag_reg.tag      = reg2hw.tag_1117.q;
  assign rcache_line[4][93].tag_reg.qe       = reg2hw.tag_1117.qe;
  assign rcache_line[4][93].tag_reg.re       = reg2hw.tag_1117.re;
  assign rcache_line[4][93].status_reg.status = reg2hw.status_1117.q;//status_reg_t'(reg2hw.status_1117.q);
  assign rcache_line[4][93].status_reg.qe    = reg2hw.status_1117.qe;
  assign rcache_line[4][93].status_reg.re    = reg2hw.status_1117.re;


  assign rcache_line[4][94].tag_reg.tag      = reg2hw.tag_1118.q;
  assign rcache_line[4][94].tag_reg.qe       = reg2hw.tag_1118.qe;
  assign rcache_line[4][94].tag_reg.re       = reg2hw.tag_1118.re;
  assign rcache_line[4][94].status_reg.status = reg2hw.status_1118.q;//status_reg_t'(reg2hw.status_1118.q);
  assign rcache_line[4][94].status_reg.qe    = reg2hw.status_1118.qe;
  assign rcache_line[4][94].status_reg.re    = reg2hw.status_1118.re;


  assign rcache_line[4][95].tag_reg.tag      = reg2hw.tag_1119.q;
  assign rcache_line[4][95].tag_reg.qe       = reg2hw.tag_1119.qe;
  assign rcache_line[4][95].tag_reg.re       = reg2hw.tag_1119.re;
  assign rcache_line[4][95].status_reg.status = reg2hw.status_1119.q;//status_reg_t'(reg2hw.status_1119.q);
  assign rcache_line[4][95].status_reg.qe    = reg2hw.status_1119.qe;
  assign rcache_line[4][95].status_reg.re    = reg2hw.status_1119.re;


  assign rcache_line[4][96].tag_reg.tag      = reg2hw.tag_1120.q;
  assign rcache_line[4][96].tag_reg.qe       = reg2hw.tag_1120.qe;
  assign rcache_line[4][96].tag_reg.re       = reg2hw.tag_1120.re;
  assign rcache_line[4][96].status_reg.status = reg2hw.status_1120.q;//status_reg_t'(reg2hw.status_1120.q);
  assign rcache_line[4][96].status_reg.qe    = reg2hw.status_1120.qe;
  assign rcache_line[4][96].status_reg.re    = reg2hw.status_1120.re;


  assign rcache_line[4][97].tag_reg.tag      = reg2hw.tag_1121.q;
  assign rcache_line[4][97].tag_reg.qe       = reg2hw.tag_1121.qe;
  assign rcache_line[4][97].tag_reg.re       = reg2hw.tag_1121.re;
  assign rcache_line[4][97].status_reg.status = reg2hw.status_1121.q;//status_reg_t'(reg2hw.status_1121.q);
  assign rcache_line[4][97].status_reg.qe    = reg2hw.status_1121.qe;
  assign rcache_line[4][97].status_reg.re    = reg2hw.status_1121.re;


  assign rcache_line[4][98].tag_reg.tag      = reg2hw.tag_1122.q;
  assign rcache_line[4][98].tag_reg.qe       = reg2hw.tag_1122.qe;
  assign rcache_line[4][98].tag_reg.re       = reg2hw.tag_1122.re;
  assign rcache_line[4][98].status_reg.status = reg2hw.status_1122.q;//status_reg_t'(reg2hw.status_1122.q);
  assign rcache_line[4][98].status_reg.qe    = reg2hw.status_1122.qe;
  assign rcache_line[4][98].status_reg.re    = reg2hw.status_1122.re;


  assign rcache_line[4][99].tag_reg.tag      = reg2hw.tag_1123.q;
  assign rcache_line[4][99].tag_reg.qe       = reg2hw.tag_1123.qe;
  assign rcache_line[4][99].tag_reg.re       = reg2hw.tag_1123.re;
  assign rcache_line[4][99].status_reg.status = reg2hw.status_1123.q;//status_reg_t'(reg2hw.status_1123.q);
  assign rcache_line[4][99].status_reg.qe    = reg2hw.status_1123.qe;
  assign rcache_line[4][99].status_reg.re    = reg2hw.status_1123.re;


  assign rcache_line[4][100].tag_reg.tag      = reg2hw.tag_1124.q;
  assign rcache_line[4][100].tag_reg.qe       = reg2hw.tag_1124.qe;
  assign rcache_line[4][100].tag_reg.re       = reg2hw.tag_1124.re;
  assign rcache_line[4][100].status_reg.status = reg2hw.status_1124.q;//status_reg_t'(reg2hw.status_1124.q);
  assign rcache_line[4][100].status_reg.qe    = reg2hw.status_1124.qe;
  assign rcache_line[4][100].status_reg.re    = reg2hw.status_1124.re;


  assign rcache_line[4][101].tag_reg.tag      = reg2hw.tag_1125.q;
  assign rcache_line[4][101].tag_reg.qe       = reg2hw.tag_1125.qe;
  assign rcache_line[4][101].tag_reg.re       = reg2hw.tag_1125.re;
  assign rcache_line[4][101].status_reg.status = reg2hw.status_1125.q;//status_reg_t'(reg2hw.status_1125.q);
  assign rcache_line[4][101].status_reg.qe    = reg2hw.status_1125.qe;
  assign rcache_line[4][101].status_reg.re    = reg2hw.status_1125.re;


  assign rcache_line[4][102].tag_reg.tag      = reg2hw.tag_1126.q;
  assign rcache_line[4][102].tag_reg.qe       = reg2hw.tag_1126.qe;
  assign rcache_line[4][102].tag_reg.re       = reg2hw.tag_1126.re;
  assign rcache_line[4][102].status_reg.status = reg2hw.status_1126.q;//status_reg_t'(reg2hw.status_1126.q);
  assign rcache_line[4][102].status_reg.qe    = reg2hw.status_1126.qe;
  assign rcache_line[4][102].status_reg.re    = reg2hw.status_1126.re;


  assign rcache_line[4][103].tag_reg.tag      = reg2hw.tag_1127.q;
  assign rcache_line[4][103].tag_reg.qe       = reg2hw.tag_1127.qe;
  assign rcache_line[4][103].tag_reg.re       = reg2hw.tag_1127.re;
  assign rcache_line[4][103].status_reg.status = reg2hw.status_1127.q;//status_reg_t'(reg2hw.status_1127.q);
  assign rcache_line[4][103].status_reg.qe    = reg2hw.status_1127.qe;
  assign rcache_line[4][103].status_reg.re    = reg2hw.status_1127.re;


  assign rcache_line[4][104].tag_reg.tag      = reg2hw.tag_1128.q;
  assign rcache_line[4][104].tag_reg.qe       = reg2hw.tag_1128.qe;
  assign rcache_line[4][104].tag_reg.re       = reg2hw.tag_1128.re;
  assign rcache_line[4][104].status_reg.status = reg2hw.status_1128.q;//status_reg_t'(reg2hw.status_1128.q);
  assign rcache_line[4][104].status_reg.qe    = reg2hw.status_1128.qe;
  assign rcache_line[4][104].status_reg.re    = reg2hw.status_1128.re;


  assign rcache_line[4][105].tag_reg.tag      = reg2hw.tag_1129.q;
  assign rcache_line[4][105].tag_reg.qe       = reg2hw.tag_1129.qe;
  assign rcache_line[4][105].tag_reg.re       = reg2hw.tag_1129.re;
  assign rcache_line[4][105].status_reg.status = reg2hw.status_1129.q;//status_reg_t'(reg2hw.status_1129.q);
  assign rcache_line[4][105].status_reg.qe    = reg2hw.status_1129.qe;
  assign rcache_line[4][105].status_reg.re    = reg2hw.status_1129.re;


  assign rcache_line[4][106].tag_reg.tag      = reg2hw.tag_1130.q;
  assign rcache_line[4][106].tag_reg.qe       = reg2hw.tag_1130.qe;
  assign rcache_line[4][106].tag_reg.re       = reg2hw.tag_1130.re;
  assign rcache_line[4][106].status_reg.status = reg2hw.status_1130.q;//status_reg_t'(reg2hw.status_1130.q);
  assign rcache_line[4][106].status_reg.qe    = reg2hw.status_1130.qe;
  assign rcache_line[4][106].status_reg.re    = reg2hw.status_1130.re;


  assign rcache_line[4][107].tag_reg.tag      = reg2hw.tag_1131.q;
  assign rcache_line[4][107].tag_reg.qe       = reg2hw.tag_1131.qe;
  assign rcache_line[4][107].tag_reg.re       = reg2hw.tag_1131.re;
  assign rcache_line[4][107].status_reg.status = reg2hw.status_1131.q;//status_reg_t'(reg2hw.status_1131.q);
  assign rcache_line[4][107].status_reg.qe    = reg2hw.status_1131.qe;
  assign rcache_line[4][107].status_reg.re    = reg2hw.status_1131.re;


  assign rcache_line[4][108].tag_reg.tag      = reg2hw.tag_1132.q;
  assign rcache_line[4][108].tag_reg.qe       = reg2hw.tag_1132.qe;
  assign rcache_line[4][108].tag_reg.re       = reg2hw.tag_1132.re;
  assign rcache_line[4][108].status_reg.status = reg2hw.status_1132.q;//status_reg_t'(reg2hw.status_1132.q);
  assign rcache_line[4][108].status_reg.qe    = reg2hw.status_1132.qe;
  assign rcache_line[4][108].status_reg.re    = reg2hw.status_1132.re;


  assign rcache_line[4][109].tag_reg.tag      = reg2hw.tag_1133.q;
  assign rcache_line[4][109].tag_reg.qe       = reg2hw.tag_1133.qe;
  assign rcache_line[4][109].tag_reg.re       = reg2hw.tag_1133.re;
  assign rcache_line[4][109].status_reg.status = reg2hw.status_1133.q;//status_reg_t'(reg2hw.status_1133.q);
  assign rcache_line[4][109].status_reg.qe    = reg2hw.status_1133.qe;
  assign rcache_line[4][109].status_reg.re    = reg2hw.status_1133.re;


  assign rcache_line[4][110].tag_reg.tag      = reg2hw.tag_1134.q;
  assign rcache_line[4][110].tag_reg.qe       = reg2hw.tag_1134.qe;
  assign rcache_line[4][110].tag_reg.re       = reg2hw.tag_1134.re;
  assign rcache_line[4][110].status_reg.status = reg2hw.status_1134.q;//status_reg_t'(reg2hw.status_1134.q);
  assign rcache_line[4][110].status_reg.qe    = reg2hw.status_1134.qe;
  assign rcache_line[4][110].status_reg.re    = reg2hw.status_1134.re;


  assign rcache_line[4][111].tag_reg.tag      = reg2hw.tag_1135.q;
  assign rcache_line[4][111].tag_reg.qe       = reg2hw.tag_1135.qe;
  assign rcache_line[4][111].tag_reg.re       = reg2hw.tag_1135.re;
  assign rcache_line[4][111].status_reg.status = reg2hw.status_1135.q;//status_reg_t'(reg2hw.status_1135.q);
  assign rcache_line[4][111].status_reg.qe    = reg2hw.status_1135.qe;
  assign rcache_line[4][111].status_reg.re    = reg2hw.status_1135.re;


  assign rcache_line[4][112].tag_reg.tag      = reg2hw.tag_1136.q;
  assign rcache_line[4][112].tag_reg.qe       = reg2hw.tag_1136.qe;
  assign rcache_line[4][112].tag_reg.re       = reg2hw.tag_1136.re;
  assign rcache_line[4][112].status_reg.status = reg2hw.status_1136.q;//status_reg_t'(reg2hw.status_1136.q);
  assign rcache_line[4][112].status_reg.qe    = reg2hw.status_1136.qe;
  assign rcache_line[4][112].status_reg.re    = reg2hw.status_1136.re;


  assign rcache_line[4][113].tag_reg.tag      = reg2hw.tag_1137.q;
  assign rcache_line[4][113].tag_reg.qe       = reg2hw.tag_1137.qe;
  assign rcache_line[4][113].tag_reg.re       = reg2hw.tag_1137.re;
  assign rcache_line[4][113].status_reg.status = reg2hw.status_1137.q;//status_reg_t'(reg2hw.status_1137.q);
  assign rcache_line[4][113].status_reg.qe    = reg2hw.status_1137.qe;
  assign rcache_line[4][113].status_reg.re    = reg2hw.status_1137.re;


  assign rcache_line[4][114].tag_reg.tag      = reg2hw.tag_1138.q;
  assign rcache_line[4][114].tag_reg.qe       = reg2hw.tag_1138.qe;
  assign rcache_line[4][114].tag_reg.re       = reg2hw.tag_1138.re;
  assign rcache_line[4][114].status_reg.status = reg2hw.status_1138.q;//status_reg_t'(reg2hw.status_1138.q);
  assign rcache_line[4][114].status_reg.qe    = reg2hw.status_1138.qe;
  assign rcache_line[4][114].status_reg.re    = reg2hw.status_1138.re;


  assign rcache_line[4][115].tag_reg.tag      = reg2hw.tag_1139.q;
  assign rcache_line[4][115].tag_reg.qe       = reg2hw.tag_1139.qe;
  assign rcache_line[4][115].tag_reg.re       = reg2hw.tag_1139.re;
  assign rcache_line[4][115].status_reg.status = reg2hw.status_1139.q;//status_reg_t'(reg2hw.status_1139.q);
  assign rcache_line[4][115].status_reg.qe    = reg2hw.status_1139.qe;
  assign rcache_line[4][115].status_reg.re    = reg2hw.status_1139.re;


  assign rcache_line[4][116].tag_reg.tag      = reg2hw.tag_1140.q;
  assign rcache_line[4][116].tag_reg.qe       = reg2hw.tag_1140.qe;
  assign rcache_line[4][116].tag_reg.re       = reg2hw.tag_1140.re;
  assign rcache_line[4][116].status_reg.status = reg2hw.status_1140.q;//status_reg_t'(reg2hw.status_1140.q);
  assign rcache_line[4][116].status_reg.qe    = reg2hw.status_1140.qe;
  assign rcache_line[4][116].status_reg.re    = reg2hw.status_1140.re;


  assign rcache_line[4][117].tag_reg.tag      = reg2hw.tag_1141.q;
  assign rcache_line[4][117].tag_reg.qe       = reg2hw.tag_1141.qe;
  assign rcache_line[4][117].tag_reg.re       = reg2hw.tag_1141.re;
  assign rcache_line[4][117].status_reg.status = reg2hw.status_1141.q;//status_reg_t'(reg2hw.status_1141.q);
  assign rcache_line[4][117].status_reg.qe    = reg2hw.status_1141.qe;
  assign rcache_line[4][117].status_reg.re    = reg2hw.status_1141.re;


  assign rcache_line[4][118].tag_reg.tag      = reg2hw.tag_1142.q;
  assign rcache_line[4][118].tag_reg.qe       = reg2hw.tag_1142.qe;
  assign rcache_line[4][118].tag_reg.re       = reg2hw.tag_1142.re;
  assign rcache_line[4][118].status_reg.status = reg2hw.status_1142.q;//status_reg_t'(reg2hw.status_1142.q);
  assign rcache_line[4][118].status_reg.qe    = reg2hw.status_1142.qe;
  assign rcache_line[4][118].status_reg.re    = reg2hw.status_1142.re;


  assign rcache_line[4][119].tag_reg.tag      = reg2hw.tag_1143.q;
  assign rcache_line[4][119].tag_reg.qe       = reg2hw.tag_1143.qe;
  assign rcache_line[4][119].tag_reg.re       = reg2hw.tag_1143.re;
  assign rcache_line[4][119].status_reg.status = reg2hw.status_1143.q;//status_reg_t'(reg2hw.status_1143.q);
  assign rcache_line[4][119].status_reg.qe    = reg2hw.status_1143.qe;
  assign rcache_line[4][119].status_reg.re    = reg2hw.status_1143.re;


  assign rcache_line[4][120].tag_reg.tag      = reg2hw.tag_1144.q;
  assign rcache_line[4][120].tag_reg.qe       = reg2hw.tag_1144.qe;
  assign rcache_line[4][120].tag_reg.re       = reg2hw.tag_1144.re;
  assign rcache_line[4][120].status_reg.status = reg2hw.status_1144.q;//status_reg_t'(reg2hw.status_1144.q);
  assign rcache_line[4][120].status_reg.qe    = reg2hw.status_1144.qe;
  assign rcache_line[4][120].status_reg.re    = reg2hw.status_1144.re;


  assign rcache_line[4][121].tag_reg.tag      = reg2hw.tag_1145.q;
  assign rcache_line[4][121].tag_reg.qe       = reg2hw.tag_1145.qe;
  assign rcache_line[4][121].tag_reg.re       = reg2hw.tag_1145.re;
  assign rcache_line[4][121].status_reg.status = reg2hw.status_1145.q;//status_reg_t'(reg2hw.status_1145.q);
  assign rcache_line[4][121].status_reg.qe    = reg2hw.status_1145.qe;
  assign rcache_line[4][121].status_reg.re    = reg2hw.status_1145.re;


  assign rcache_line[4][122].tag_reg.tag      = reg2hw.tag_1146.q;
  assign rcache_line[4][122].tag_reg.qe       = reg2hw.tag_1146.qe;
  assign rcache_line[4][122].tag_reg.re       = reg2hw.tag_1146.re;
  assign rcache_line[4][122].status_reg.status = reg2hw.status_1146.q;//status_reg_t'(reg2hw.status_1146.q);
  assign rcache_line[4][122].status_reg.qe    = reg2hw.status_1146.qe;
  assign rcache_line[4][122].status_reg.re    = reg2hw.status_1146.re;


  assign rcache_line[4][123].tag_reg.tag      = reg2hw.tag_1147.q;
  assign rcache_line[4][123].tag_reg.qe       = reg2hw.tag_1147.qe;
  assign rcache_line[4][123].tag_reg.re       = reg2hw.tag_1147.re;
  assign rcache_line[4][123].status_reg.status = reg2hw.status_1147.q;//status_reg_t'(reg2hw.status_1147.q);
  assign rcache_line[4][123].status_reg.qe    = reg2hw.status_1147.qe;
  assign rcache_line[4][123].status_reg.re    = reg2hw.status_1147.re;


  assign rcache_line[4][124].tag_reg.tag      = reg2hw.tag_1148.q;
  assign rcache_line[4][124].tag_reg.qe       = reg2hw.tag_1148.qe;
  assign rcache_line[4][124].tag_reg.re       = reg2hw.tag_1148.re;
  assign rcache_line[4][124].status_reg.status = reg2hw.status_1148.q;//status_reg_t'(reg2hw.status_1148.q);
  assign rcache_line[4][124].status_reg.qe    = reg2hw.status_1148.qe;
  assign rcache_line[4][124].status_reg.re    = reg2hw.status_1148.re;


  assign rcache_line[4][125].tag_reg.tag      = reg2hw.tag_1149.q;
  assign rcache_line[4][125].tag_reg.qe       = reg2hw.tag_1149.qe;
  assign rcache_line[4][125].tag_reg.re       = reg2hw.tag_1149.re;
  assign rcache_line[4][125].status_reg.status = reg2hw.status_1149.q;//status_reg_t'(reg2hw.status_1149.q);
  assign rcache_line[4][125].status_reg.qe    = reg2hw.status_1149.qe;
  assign rcache_line[4][125].status_reg.re    = reg2hw.status_1149.re;


  assign rcache_line[4][126].tag_reg.tag      = reg2hw.tag_1150.q;
  assign rcache_line[4][126].tag_reg.qe       = reg2hw.tag_1150.qe;
  assign rcache_line[4][126].tag_reg.re       = reg2hw.tag_1150.re;
  assign rcache_line[4][126].status_reg.status = reg2hw.status_1150.q;//status_reg_t'(reg2hw.status_1150.q);
  assign rcache_line[4][126].status_reg.qe    = reg2hw.status_1150.qe;
  assign rcache_line[4][126].status_reg.re    = reg2hw.status_1150.re;


  assign rcache_line[4][127].tag_reg.tag      = reg2hw.tag_1151.q;
  assign rcache_line[4][127].tag_reg.qe       = reg2hw.tag_1151.qe;
  assign rcache_line[4][127].tag_reg.re       = reg2hw.tag_1151.re;
  assign rcache_line[4][127].status_reg.status = reg2hw.status_1151.q;//status_reg_t'(reg2hw.status_1151.q);
  assign rcache_line[4][127].status_reg.qe    = reg2hw.status_1151.qe;
  assign rcache_line[4][127].status_reg.re    = reg2hw.status_1151.re;


  assign rcache_line[4][128].tag_reg.tag      = reg2hw.tag_1152.q;
  assign rcache_line[4][128].tag_reg.qe       = reg2hw.tag_1152.qe;
  assign rcache_line[4][128].tag_reg.re       = reg2hw.tag_1152.re;
  assign rcache_line[4][128].status_reg.status = reg2hw.status_1152.q;//status_reg_t'(reg2hw.status_1152.q);
  assign rcache_line[4][128].status_reg.qe    = reg2hw.status_1152.qe;
  assign rcache_line[4][128].status_reg.re    = reg2hw.status_1152.re;


  assign rcache_line[4][129].tag_reg.tag      = reg2hw.tag_1153.q;
  assign rcache_line[4][129].tag_reg.qe       = reg2hw.tag_1153.qe;
  assign rcache_line[4][129].tag_reg.re       = reg2hw.tag_1153.re;
  assign rcache_line[4][129].status_reg.status = reg2hw.status_1153.q;//status_reg_t'(reg2hw.status_1153.q);
  assign rcache_line[4][129].status_reg.qe    = reg2hw.status_1153.qe;
  assign rcache_line[4][129].status_reg.re    = reg2hw.status_1153.re;


  assign rcache_line[4][130].tag_reg.tag      = reg2hw.tag_1154.q;
  assign rcache_line[4][130].tag_reg.qe       = reg2hw.tag_1154.qe;
  assign rcache_line[4][130].tag_reg.re       = reg2hw.tag_1154.re;
  assign rcache_line[4][130].status_reg.status = reg2hw.status_1154.q;//status_reg_t'(reg2hw.status_1154.q);
  assign rcache_line[4][130].status_reg.qe    = reg2hw.status_1154.qe;
  assign rcache_line[4][130].status_reg.re    = reg2hw.status_1154.re;


  assign rcache_line[4][131].tag_reg.tag      = reg2hw.tag_1155.q;
  assign rcache_line[4][131].tag_reg.qe       = reg2hw.tag_1155.qe;
  assign rcache_line[4][131].tag_reg.re       = reg2hw.tag_1155.re;
  assign rcache_line[4][131].status_reg.status = reg2hw.status_1155.q;//status_reg_t'(reg2hw.status_1155.q);
  assign rcache_line[4][131].status_reg.qe    = reg2hw.status_1155.qe;
  assign rcache_line[4][131].status_reg.re    = reg2hw.status_1155.re;


  assign rcache_line[4][132].tag_reg.tag      = reg2hw.tag_1156.q;
  assign rcache_line[4][132].tag_reg.qe       = reg2hw.tag_1156.qe;
  assign rcache_line[4][132].tag_reg.re       = reg2hw.tag_1156.re;
  assign rcache_line[4][132].status_reg.status = reg2hw.status_1156.q;//status_reg_t'(reg2hw.status_1156.q);
  assign rcache_line[4][132].status_reg.qe    = reg2hw.status_1156.qe;
  assign rcache_line[4][132].status_reg.re    = reg2hw.status_1156.re;


  assign rcache_line[4][133].tag_reg.tag      = reg2hw.tag_1157.q;
  assign rcache_line[4][133].tag_reg.qe       = reg2hw.tag_1157.qe;
  assign rcache_line[4][133].tag_reg.re       = reg2hw.tag_1157.re;
  assign rcache_line[4][133].status_reg.status = reg2hw.status_1157.q;//status_reg_t'(reg2hw.status_1157.q);
  assign rcache_line[4][133].status_reg.qe    = reg2hw.status_1157.qe;
  assign rcache_line[4][133].status_reg.re    = reg2hw.status_1157.re;


  assign rcache_line[4][134].tag_reg.tag      = reg2hw.tag_1158.q;
  assign rcache_line[4][134].tag_reg.qe       = reg2hw.tag_1158.qe;
  assign rcache_line[4][134].tag_reg.re       = reg2hw.tag_1158.re;
  assign rcache_line[4][134].status_reg.status = reg2hw.status_1158.q;//status_reg_t'(reg2hw.status_1158.q);
  assign rcache_line[4][134].status_reg.qe    = reg2hw.status_1158.qe;
  assign rcache_line[4][134].status_reg.re    = reg2hw.status_1158.re;


  assign rcache_line[4][135].tag_reg.tag      = reg2hw.tag_1159.q;
  assign rcache_line[4][135].tag_reg.qe       = reg2hw.tag_1159.qe;
  assign rcache_line[4][135].tag_reg.re       = reg2hw.tag_1159.re;
  assign rcache_line[4][135].status_reg.status = reg2hw.status_1159.q;//status_reg_t'(reg2hw.status_1159.q);
  assign rcache_line[4][135].status_reg.qe    = reg2hw.status_1159.qe;
  assign rcache_line[4][135].status_reg.re    = reg2hw.status_1159.re;


  assign rcache_line[4][136].tag_reg.tag      = reg2hw.tag_1160.q;
  assign rcache_line[4][136].tag_reg.qe       = reg2hw.tag_1160.qe;
  assign rcache_line[4][136].tag_reg.re       = reg2hw.tag_1160.re;
  assign rcache_line[4][136].status_reg.status = reg2hw.status_1160.q;//status_reg_t'(reg2hw.status_1160.q);
  assign rcache_line[4][136].status_reg.qe    = reg2hw.status_1160.qe;
  assign rcache_line[4][136].status_reg.re    = reg2hw.status_1160.re;


  assign rcache_line[4][137].tag_reg.tag      = reg2hw.tag_1161.q;
  assign rcache_line[4][137].tag_reg.qe       = reg2hw.tag_1161.qe;
  assign rcache_line[4][137].tag_reg.re       = reg2hw.tag_1161.re;
  assign rcache_line[4][137].status_reg.status = reg2hw.status_1161.q;//status_reg_t'(reg2hw.status_1161.q);
  assign rcache_line[4][137].status_reg.qe    = reg2hw.status_1161.qe;
  assign rcache_line[4][137].status_reg.re    = reg2hw.status_1161.re;


  assign rcache_line[4][138].tag_reg.tag      = reg2hw.tag_1162.q;
  assign rcache_line[4][138].tag_reg.qe       = reg2hw.tag_1162.qe;
  assign rcache_line[4][138].tag_reg.re       = reg2hw.tag_1162.re;
  assign rcache_line[4][138].status_reg.status = reg2hw.status_1162.q;//status_reg_t'(reg2hw.status_1162.q);
  assign rcache_line[4][138].status_reg.qe    = reg2hw.status_1162.qe;
  assign rcache_line[4][138].status_reg.re    = reg2hw.status_1162.re;


  assign rcache_line[4][139].tag_reg.tag      = reg2hw.tag_1163.q;
  assign rcache_line[4][139].tag_reg.qe       = reg2hw.tag_1163.qe;
  assign rcache_line[4][139].tag_reg.re       = reg2hw.tag_1163.re;
  assign rcache_line[4][139].status_reg.status = reg2hw.status_1163.q;//status_reg_t'(reg2hw.status_1163.q);
  assign rcache_line[4][139].status_reg.qe    = reg2hw.status_1163.qe;
  assign rcache_line[4][139].status_reg.re    = reg2hw.status_1163.re;


  assign rcache_line[4][140].tag_reg.tag      = reg2hw.tag_1164.q;
  assign rcache_line[4][140].tag_reg.qe       = reg2hw.tag_1164.qe;
  assign rcache_line[4][140].tag_reg.re       = reg2hw.tag_1164.re;
  assign rcache_line[4][140].status_reg.status = reg2hw.status_1164.q;//status_reg_t'(reg2hw.status_1164.q);
  assign rcache_line[4][140].status_reg.qe    = reg2hw.status_1164.qe;
  assign rcache_line[4][140].status_reg.re    = reg2hw.status_1164.re;


  assign rcache_line[4][141].tag_reg.tag      = reg2hw.tag_1165.q;
  assign rcache_line[4][141].tag_reg.qe       = reg2hw.tag_1165.qe;
  assign rcache_line[4][141].tag_reg.re       = reg2hw.tag_1165.re;
  assign rcache_line[4][141].status_reg.status = reg2hw.status_1165.q;//status_reg_t'(reg2hw.status_1165.q);
  assign rcache_line[4][141].status_reg.qe    = reg2hw.status_1165.qe;
  assign rcache_line[4][141].status_reg.re    = reg2hw.status_1165.re;


  assign rcache_line[4][142].tag_reg.tag      = reg2hw.tag_1166.q;
  assign rcache_line[4][142].tag_reg.qe       = reg2hw.tag_1166.qe;
  assign rcache_line[4][142].tag_reg.re       = reg2hw.tag_1166.re;
  assign rcache_line[4][142].status_reg.status = reg2hw.status_1166.q;//status_reg_t'(reg2hw.status_1166.q);
  assign rcache_line[4][142].status_reg.qe    = reg2hw.status_1166.qe;
  assign rcache_line[4][142].status_reg.re    = reg2hw.status_1166.re;


  assign rcache_line[4][143].tag_reg.tag      = reg2hw.tag_1167.q;
  assign rcache_line[4][143].tag_reg.qe       = reg2hw.tag_1167.qe;
  assign rcache_line[4][143].tag_reg.re       = reg2hw.tag_1167.re;
  assign rcache_line[4][143].status_reg.status = reg2hw.status_1167.q;//status_reg_t'(reg2hw.status_1167.q);
  assign rcache_line[4][143].status_reg.qe    = reg2hw.status_1167.qe;
  assign rcache_line[4][143].status_reg.re    = reg2hw.status_1167.re;


  assign rcache_line[4][144].tag_reg.tag      = reg2hw.tag_1168.q;
  assign rcache_line[4][144].tag_reg.qe       = reg2hw.tag_1168.qe;
  assign rcache_line[4][144].tag_reg.re       = reg2hw.tag_1168.re;
  assign rcache_line[4][144].status_reg.status = reg2hw.status_1168.q;//status_reg_t'(reg2hw.status_1168.q);
  assign rcache_line[4][144].status_reg.qe    = reg2hw.status_1168.qe;
  assign rcache_line[4][144].status_reg.re    = reg2hw.status_1168.re;


  assign rcache_line[4][145].tag_reg.tag      = reg2hw.tag_1169.q;
  assign rcache_line[4][145].tag_reg.qe       = reg2hw.tag_1169.qe;
  assign rcache_line[4][145].tag_reg.re       = reg2hw.tag_1169.re;
  assign rcache_line[4][145].status_reg.status = reg2hw.status_1169.q;//status_reg_t'(reg2hw.status_1169.q);
  assign rcache_line[4][145].status_reg.qe    = reg2hw.status_1169.qe;
  assign rcache_line[4][145].status_reg.re    = reg2hw.status_1169.re;


  assign rcache_line[4][146].tag_reg.tag      = reg2hw.tag_1170.q;
  assign rcache_line[4][146].tag_reg.qe       = reg2hw.tag_1170.qe;
  assign rcache_line[4][146].tag_reg.re       = reg2hw.tag_1170.re;
  assign rcache_line[4][146].status_reg.status = reg2hw.status_1170.q;//status_reg_t'(reg2hw.status_1170.q);
  assign rcache_line[4][146].status_reg.qe    = reg2hw.status_1170.qe;
  assign rcache_line[4][146].status_reg.re    = reg2hw.status_1170.re;


  assign rcache_line[4][147].tag_reg.tag      = reg2hw.tag_1171.q;
  assign rcache_line[4][147].tag_reg.qe       = reg2hw.tag_1171.qe;
  assign rcache_line[4][147].tag_reg.re       = reg2hw.tag_1171.re;
  assign rcache_line[4][147].status_reg.status = reg2hw.status_1171.q;//status_reg_t'(reg2hw.status_1171.q);
  assign rcache_line[4][147].status_reg.qe    = reg2hw.status_1171.qe;
  assign rcache_line[4][147].status_reg.re    = reg2hw.status_1171.re;


  assign rcache_line[4][148].tag_reg.tag      = reg2hw.tag_1172.q;
  assign rcache_line[4][148].tag_reg.qe       = reg2hw.tag_1172.qe;
  assign rcache_line[4][148].tag_reg.re       = reg2hw.tag_1172.re;
  assign rcache_line[4][148].status_reg.status = reg2hw.status_1172.q;//status_reg_t'(reg2hw.status_1172.q);
  assign rcache_line[4][148].status_reg.qe    = reg2hw.status_1172.qe;
  assign rcache_line[4][148].status_reg.re    = reg2hw.status_1172.re;


  assign rcache_line[4][149].tag_reg.tag      = reg2hw.tag_1173.q;
  assign rcache_line[4][149].tag_reg.qe       = reg2hw.tag_1173.qe;
  assign rcache_line[4][149].tag_reg.re       = reg2hw.tag_1173.re;
  assign rcache_line[4][149].status_reg.status = reg2hw.status_1173.q;//status_reg_t'(reg2hw.status_1173.q);
  assign rcache_line[4][149].status_reg.qe    = reg2hw.status_1173.qe;
  assign rcache_line[4][149].status_reg.re    = reg2hw.status_1173.re;


  assign rcache_line[4][150].tag_reg.tag      = reg2hw.tag_1174.q;
  assign rcache_line[4][150].tag_reg.qe       = reg2hw.tag_1174.qe;
  assign rcache_line[4][150].tag_reg.re       = reg2hw.tag_1174.re;
  assign rcache_line[4][150].status_reg.status = reg2hw.status_1174.q;//status_reg_t'(reg2hw.status_1174.q);
  assign rcache_line[4][150].status_reg.qe    = reg2hw.status_1174.qe;
  assign rcache_line[4][150].status_reg.re    = reg2hw.status_1174.re;


  assign rcache_line[4][151].tag_reg.tag      = reg2hw.tag_1175.q;
  assign rcache_line[4][151].tag_reg.qe       = reg2hw.tag_1175.qe;
  assign rcache_line[4][151].tag_reg.re       = reg2hw.tag_1175.re;
  assign rcache_line[4][151].status_reg.status = reg2hw.status_1175.q;//status_reg_t'(reg2hw.status_1175.q);
  assign rcache_line[4][151].status_reg.qe    = reg2hw.status_1175.qe;
  assign rcache_line[4][151].status_reg.re    = reg2hw.status_1175.re;


  assign rcache_line[4][152].tag_reg.tag      = reg2hw.tag_1176.q;
  assign rcache_line[4][152].tag_reg.qe       = reg2hw.tag_1176.qe;
  assign rcache_line[4][152].tag_reg.re       = reg2hw.tag_1176.re;
  assign rcache_line[4][152].status_reg.status = reg2hw.status_1176.q;//status_reg_t'(reg2hw.status_1176.q);
  assign rcache_line[4][152].status_reg.qe    = reg2hw.status_1176.qe;
  assign rcache_line[4][152].status_reg.re    = reg2hw.status_1176.re;


  assign rcache_line[4][153].tag_reg.tag      = reg2hw.tag_1177.q;
  assign rcache_line[4][153].tag_reg.qe       = reg2hw.tag_1177.qe;
  assign rcache_line[4][153].tag_reg.re       = reg2hw.tag_1177.re;
  assign rcache_line[4][153].status_reg.status = reg2hw.status_1177.q;//status_reg_t'(reg2hw.status_1177.q);
  assign rcache_line[4][153].status_reg.qe    = reg2hw.status_1177.qe;
  assign rcache_line[4][153].status_reg.re    = reg2hw.status_1177.re;


  assign rcache_line[4][154].tag_reg.tag      = reg2hw.tag_1178.q;
  assign rcache_line[4][154].tag_reg.qe       = reg2hw.tag_1178.qe;
  assign rcache_line[4][154].tag_reg.re       = reg2hw.tag_1178.re;
  assign rcache_line[4][154].status_reg.status = reg2hw.status_1178.q;//status_reg_t'(reg2hw.status_1178.q);
  assign rcache_line[4][154].status_reg.qe    = reg2hw.status_1178.qe;
  assign rcache_line[4][154].status_reg.re    = reg2hw.status_1178.re;


  assign rcache_line[4][155].tag_reg.tag      = reg2hw.tag_1179.q;
  assign rcache_line[4][155].tag_reg.qe       = reg2hw.tag_1179.qe;
  assign rcache_line[4][155].tag_reg.re       = reg2hw.tag_1179.re;
  assign rcache_line[4][155].status_reg.status = reg2hw.status_1179.q;//status_reg_t'(reg2hw.status_1179.q);
  assign rcache_line[4][155].status_reg.qe    = reg2hw.status_1179.qe;
  assign rcache_line[4][155].status_reg.re    = reg2hw.status_1179.re;


  assign rcache_line[4][156].tag_reg.tag      = reg2hw.tag_1180.q;
  assign rcache_line[4][156].tag_reg.qe       = reg2hw.tag_1180.qe;
  assign rcache_line[4][156].tag_reg.re       = reg2hw.tag_1180.re;
  assign rcache_line[4][156].status_reg.status = reg2hw.status_1180.q;//status_reg_t'(reg2hw.status_1180.q);
  assign rcache_line[4][156].status_reg.qe    = reg2hw.status_1180.qe;
  assign rcache_line[4][156].status_reg.re    = reg2hw.status_1180.re;


  assign rcache_line[4][157].tag_reg.tag      = reg2hw.tag_1181.q;
  assign rcache_line[4][157].tag_reg.qe       = reg2hw.tag_1181.qe;
  assign rcache_line[4][157].tag_reg.re       = reg2hw.tag_1181.re;
  assign rcache_line[4][157].status_reg.status = reg2hw.status_1181.q;//status_reg_t'(reg2hw.status_1181.q);
  assign rcache_line[4][157].status_reg.qe    = reg2hw.status_1181.qe;
  assign rcache_line[4][157].status_reg.re    = reg2hw.status_1181.re;


  assign rcache_line[4][158].tag_reg.tag      = reg2hw.tag_1182.q;
  assign rcache_line[4][158].tag_reg.qe       = reg2hw.tag_1182.qe;
  assign rcache_line[4][158].tag_reg.re       = reg2hw.tag_1182.re;
  assign rcache_line[4][158].status_reg.status = reg2hw.status_1182.q;//status_reg_t'(reg2hw.status_1182.q);
  assign rcache_line[4][158].status_reg.qe    = reg2hw.status_1182.qe;
  assign rcache_line[4][158].status_reg.re    = reg2hw.status_1182.re;


  assign rcache_line[4][159].tag_reg.tag      = reg2hw.tag_1183.q;
  assign rcache_line[4][159].tag_reg.qe       = reg2hw.tag_1183.qe;
  assign rcache_line[4][159].tag_reg.re       = reg2hw.tag_1183.re;
  assign rcache_line[4][159].status_reg.status = reg2hw.status_1183.q;//status_reg_t'(reg2hw.status_1183.q);
  assign rcache_line[4][159].status_reg.qe    = reg2hw.status_1183.qe;
  assign rcache_line[4][159].status_reg.re    = reg2hw.status_1183.re;


  assign rcache_line[4][160].tag_reg.tag      = reg2hw.tag_1184.q;
  assign rcache_line[4][160].tag_reg.qe       = reg2hw.tag_1184.qe;
  assign rcache_line[4][160].tag_reg.re       = reg2hw.tag_1184.re;
  assign rcache_line[4][160].status_reg.status = reg2hw.status_1184.q;//status_reg_t'(reg2hw.status_1184.q);
  assign rcache_line[4][160].status_reg.qe    = reg2hw.status_1184.qe;
  assign rcache_line[4][160].status_reg.re    = reg2hw.status_1184.re;


  assign rcache_line[4][161].tag_reg.tag      = reg2hw.tag_1185.q;
  assign rcache_line[4][161].tag_reg.qe       = reg2hw.tag_1185.qe;
  assign rcache_line[4][161].tag_reg.re       = reg2hw.tag_1185.re;
  assign rcache_line[4][161].status_reg.status = reg2hw.status_1185.q;//status_reg_t'(reg2hw.status_1185.q);
  assign rcache_line[4][161].status_reg.qe    = reg2hw.status_1185.qe;
  assign rcache_line[4][161].status_reg.re    = reg2hw.status_1185.re;


  assign rcache_line[4][162].tag_reg.tag      = reg2hw.tag_1186.q;
  assign rcache_line[4][162].tag_reg.qe       = reg2hw.tag_1186.qe;
  assign rcache_line[4][162].tag_reg.re       = reg2hw.tag_1186.re;
  assign rcache_line[4][162].status_reg.status = reg2hw.status_1186.q;//status_reg_t'(reg2hw.status_1186.q);
  assign rcache_line[4][162].status_reg.qe    = reg2hw.status_1186.qe;
  assign rcache_line[4][162].status_reg.re    = reg2hw.status_1186.re;


  assign rcache_line[4][163].tag_reg.tag      = reg2hw.tag_1187.q;
  assign rcache_line[4][163].tag_reg.qe       = reg2hw.tag_1187.qe;
  assign rcache_line[4][163].tag_reg.re       = reg2hw.tag_1187.re;
  assign rcache_line[4][163].status_reg.status = reg2hw.status_1187.q;//status_reg_t'(reg2hw.status_1187.q);
  assign rcache_line[4][163].status_reg.qe    = reg2hw.status_1187.qe;
  assign rcache_line[4][163].status_reg.re    = reg2hw.status_1187.re;


  assign rcache_line[4][164].tag_reg.tag      = reg2hw.tag_1188.q;
  assign rcache_line[4][164].tag_reg.qe       = reg2hw.tag_1188.qe;
  assign rcache_line[4][164].tag_reg.re       = reg2hw.tag_1188.re;
  assign rcache_line[4][164].status_reg.status = reg2hw.status_1188.q;//status_reg_t'(reg2hw.status_1188.q);
  assign rcache_line[4][164].status_reg.qe    = reg2hw.status_1188.qe;
  assign rcache_line[4][164].status_reg.re    = reg2hw.status_1188.re;


  assign rcache_line[4][165].tag_reg.tag      = reg2hw.tag_1189.q;
  assign rcache_line[4][165].tag_reg.qe       = reg2hw.tag_1189.qe;
  assign rcache_line[4][165].tag_reg.re       = reg2hw.tag_1189.re;
  assign rcache_line[4][165].status_reg.status = reg2hw.status_1189.q;//status_reg_t'(reg2hw.status_1189.q);
  assign rcache_line[4][165].status_reg.qe    = reg2hw.status_1189.qe;
  assign rcache_line[4][165].status_reg.re    = reg2hw.status_1189.re;


  assign rcache_line[4][166].tag_reg.tag      = reg2hw.tag_1190.q;
  assign rcache_line[4][166].tag_reg.qe       = reg2hw.tag_1190.qe;
  assign rcache_line[4][166].tag_reg.re       = reg2hw.tag_1190.re;
  assign rcache_line[4][166].status_reg.status = reg2hw.status_1190.q;//status_reg_t'(reg2hw.status_1190.q);
  assign rcache_line[4][166].status_reg.qe    = reg2hw.status_1190.qe;
  assign rcache_line[4][166].status_reg.re    = reg2hw.status_1190.re;


  assign rcache_line[4][167].tag_reg.tag      = reg2hw.tag_1191.q;
  assign rcache_line[4][167].tag_reg.qe       = reg2hw.tag_1191.qe;
  assign rcache_line[4][167].tag_reg.re       = reg2hw.tag_1191.re;
  assign rcache_line[4][167].status_reg.status = reg2hw.status_1191.q;//status_reg_t'(reg2hw.status_1191.q);
  assign rcache_line[4][167].status_reg.qe    = reg2hw.status_1191.qe;
  assign rcache_line[4][167].status_reg.re    = reg2hw.status_1191.re;


  assign rcache_line[4][168].tag_reg.tag      = reg2hw.tag_1192.q;
  assign rcache_line[4][168].tag_reg.qe       = reg2hw.tag_1192.qe;
  assign rcache_line[4][168].tag_reg.re       = reg2hw.tag_1192.re;
  assign rcache_line[4][168].status_reg.status = reg2hw.status_1192.q;//status_reg_t'(reg2hw.status_1192.q);
  assign rcache_line[4][168].status_reg.qe    = reg2hw.status_1192.qe;
  assign rcache_line[4][168].status_reg.re    = reg2hw.status_1192.re;


  assign rcache_line[4][169].tag_reg.tag      = reg2hw.tag_1193.q;
  assign rcache_line[4][169].tag_reg.qe       = reg2hw.tag_1193.qe;
  assign rcache_line[4][169].tag_reg.re       = reg2hw.tag_1193.re;
  assign rcache_line[4][169].status_reg.status = reg2hw.status_1193.q;//status_reg_t'(reg2hw.status_1193.q);
  assign rcache_line[4][169].status_reg.qe    = reg2hw.status_1193.qe;
  assign rcache_line[4][169].status_reg.re    = reg2hw.status_1193.re;


  assign rcache_line[4][170].tag_reg.tag      = reg2hw.tag_1194.q;
  assign rcache_line[4][170].tag_reg.qe       = reg2hw.tag_1194.qe;
  assign rcache_line[4][170].tag_reg.re       = reg2hw.tag_1194.re;
  assign rcache_line[4][170].status_reg.status = reg2hw.status_1194.q;//status_reg_t'(reg2hw.status_1194.q);
  assign rcache_line[4][170].status_reg.qe    = reg2hw.status_1194.qe;
  assign rcache_line[4][170].status_reg.re    = reg2hw.status_1194.re;


  assign rcache_line[4][171].tag_reg.tag      = reg2hw.tag_1195.q;
  assign rcache_line[4][171].tag_reg.qe       = reg2hw.tag_1195.qe;
  assign rcache_line[4][171].tag_reg.re       = reg2hw.tag_1195.re;
  assign rcache_line[4][171].status_reg.status = reg2hw.status_1195.q;//status_reg_t'(reg2hw.status_1195.q);
  assign rcache_line[4][171].status_reg.qe    = reg2hw.status_1195.qe;
  assign rcache_line[4][171].status_reg.re    = reg2hw.status_1195.re;


  assign rcache_line[4][172].tag_reg.tag      = reg2hw.tag_1196.q;
  assign rcache_line[4][172].tag_reg.qe       = reg2hw.tag_1196.qe;
  assign rcache_line[4][172].tag_reg.re       = reg2hw.tag_1196.re;
  assign rcache_line[4][172].status_reg.status = reg2hw.status_1196.q;//status_reg_t'(reg2hw.status_1196.q);
  assign rcache_line[4][172].status_reg.qe    = reg2hw.status_1196.qe;
  assign rcache_line[4][172].status_reg.re    = reg2hw.status_1196.re;


  assign rcache_line[4][173].tag_reg.tag      = reg2hw.tag_1197.q;
  assign rcache_line[4][173].tag_reg.qe       = reg2hw.tag_1197.qe;
  assign rcache_line[4][173].tag_reg.re       = reg2hw.tag_1197.re;
  assign rcache_line[4][173].status_reg.status = reg2hw.status_1197.q;//status_reg_t'(reg2hw.status_1197.q);
  assign rcache_line[4][173].status_reg.qe    = reg2hw.status_1197.qe;
  assign rcache_line[4][173].status_reg.re    = reg2hw.status_1197.re;


  assign rcache_line[4][174].tag_reg.tag      = reg2hw.tag_1198.q;
  assign rcache_line[4][174].tag_reg.qe       = reg2hw.tag_1198.qe;
  assign rcache_line[4][174].tag_reg.re       = reg2hw.tag_1198.re;
  assign rcache_line[4][174].status_reg.status = reg2hw.status_1198.q;//status_reg_t'(reg2hw.status_1198.q);
  assign rcache_line[4][174].status_reg.qe    = reg2hw.status_1198.qe;
  assign rcache_line[4][174].status_reg.re    = reg2hw.status_1198.re;


  assign rcache_line[4][175].tag_reg.tag      = reg2hw.tag_1199.q;
  assign rcache_line[4][175].tag_reg.qe       = reg2hw.tag_1199.qe;
  assign rcache_line[4][175].tag_reg.re       = reg2hw.tag_1199.re;
  assign rcache_line[4][175].status_reg.status = reg2hw.status_1199.q;//status_reg_t'(reg2hw.status_1199.q);
  assign rcache_line[4][175].status_reg.qe    = reg2hw.status_1199.qe;
  assign rcache_line[4][175].status_reg.re    = reg2hw.status_1199.re;


  assign rcache_line[4][176].tag_reg.tag      = reg2hw.tag_1200.q;
  assign rcache_line[4][176].tag_reg.qe       = reg2hw.tag_1200.qe;
  assign rcache_line[4][176].tag_reg.re       = reg2hw.tag_1200.re;
  assign rcache_line[4][176].status_reg.status = reg2hw.status_1200.q;//status_reg_t'(reg2hw.status_1200.q);
  assign rcache_line[4][176].status_reg.qe    = reg2hw.status_1200.qe;
  assign rcache_line[4][176].status_reg.re    = reg2hw.status_1200.re;


  assign rcache_line[4][177].tag_reg.tag      = reg2hw.tag_1201.q;
  assign rcache_line[4][177].tag_reg.qe       = reg2hw.tag_1201.qe;
  assign rcache_line[4][177].tag_reg.re       = reg2hw.tag_1201.re;
  assign rcache_line[4][177].status_reg.status = reg2hw.status_1201.q;//status_reg_t'(reg2hw.status_1201.q);
  assign rcache_line[4][177].status_reg.qe    = reg2hw.status_1201.qe;
  assign rcache_line[4][177].status_reg.re    = reg2hw.status_1201.re;


  assign rcache_line[4][178].tag_reg.tag      = reg2hw.tag_1202.q;
  assign rcache_line[4][178].tag_reg.qe       = reg2hw.tag_1202.qe;
  assign rcache_line[4][178].tag_reg.re       = reg2hw.tag_1202.re;
  assign rcache_line[4][178].status_reg.status = reg2hw.status_1202.q;//status_reg_t'(reg2hw.status_1202.q);
  assign rcache_line[4][178].status_reg.qe    = reg2hw.status_1202.qe;
  assign rcache_line[4][178].status_reg.re    = reg2hw.status_1202.re;


  assign rcache_line[4][179].tag_reg.tag      = reg2hw.tag_1203.q;
  assign rcache_line[4][179].tag_reg.qe       = reg2hw.tag_1203.qe;
  assign rcache_line[4][179].tag_reg.re       = reg2hw.tag_1203.re;
  assign rcache_line[4][179].status_reg.status = reg2hw.status_1203.q;//status_reg_t'(reg2hw.status_1203.q);
  assign rcache_line[4][179].status_reg.qe    = reg2hw.status_1203.qe;
  assign rcache_line[4][179].status_reg.re    = reg2hw.status_1203.re;


  assign rcache_line[4][180].tag_reg.tag      = reg2hw.tag_1204.q;
  assign rcache_line[4][180].tag_reg.qe       = reg2hw.tag_1204.qe;
  assign rcache_line[4][180].tag_reg.re       = reg2hw.tag_1204.re;
  assign rcache_line[4][180].status_reg.status = reg2hw.status_1204.q;//status_reg_t'(reg2hw.status_1204.q);
  assign rcache_line[4][180].status_reg.qe    = reg2hw.status_1204.qe;
  assign rcache_line[4][180].status_reg.re    = reg2hw.status_1204.re;


  assign rcache_line[4][181].tag_reg.tag      = reg2hw.tag_1205.q;
  assign rcache_line[4][181].tag_reg.qe       = reg2hw.tag_1205.qe;
  assign rcache_line[4][181].tag_reg.re       = reg2hw.tag_1205.re;
  assign rcache_line[4][181].status_reg.status = reg2hw.status_1205.q;//status_reg_t'(reg2hw.status_1205.q);
  assign rcache_line[4][181].status_reg.qe    = reg2hw.status_1205.qe;
  assign rcache_line[4][181].status_reg.re    = reg2hw.status_1205.re;


  assign rcache_line[4][182].tag_reg.tag      = reg2hw.tag_1206.q;
  assign rcache_line[4][182].tag_reg.qe       = reg2hw.tag_1206.qe;
  assign rcache_line[4][182].tag_reg.re       = reg2hw.tag_1206.re;
  assign rcache_line[4][182].status_reg.status = reg2hw.status_1206.q;//status_reg_t'(reg2hw.status_1206.q);
  assign rcache_line[4][182].status_reg.qe    = reg2hw.status_1206.qe;
  assign rcache_line[4][182].status_reg.re    = reg2hw.status_1206.re;


  assign rcache_line[4][183].tag_reg.tag      = reg2hw.tag_1207.q;
  assign rcache_line[4][183].tag_reg.qe       = reg2hw.tag_1207.qe;
  assign rcache_line[4][183].tag_reg.re       = reg2hw.tag_1207.re;
  assign rcache_line[4][183].status_reg.status = reg2hw.status_1207.q;//status_reg_t'(reg2hw.status_1207.q);
  assign rcache_line[4][183].status_reg.qe    = reg2hw.status_1207.qe;
  assign rcache_line[4][183].status_reg.re    = reg2hw.status_1207.re;


  assign rcache_line[4][184].tag_reg.tag      = reg2hw.tag_1208.q;
  assign rcache_line[4][184].tag_reg.qe       = reg2hw.tag_1208.qe;
  assign rcache_line[4][184].tag_reg.re       = reg2hw.tag_1208.re;
  assign rcache_line[4][184].status_reg.status = reg2hw.status_1208.q;//status_reg_t'(reg2hw.status_1208.q);
  assign rcache_line[4][184].status_reg.qe    = reg2hw.status_1208.qe;
  assign rcache_line[4][184].status_reg.re    = reg2hw.status_1208.re;


  assign rcache_line[4][185].tag_reg.tag      = reg2hw.tag_1209.q;
  assign rcache_line[4][185].tag_reg.qe       = reg2hw.tag_1209.qe;
  assign rcache_line[4][185].tag_reg.re       = reg2hw.tag_1209.re;
  assign rcache_line[4][185].status_reg.status = reg2hw.status_1209.q;//status_reg_t'(reg2hw.status_1209.q);
  assign rcache_line[4][185].status_reg.qe    = reg2hw.status_1209.qe;
  assign rcache_line[4][185].status_reg.re    = reg2hw.status_1209.re;


  assign rcache_line[4][186].tag_reg.tag      = reg2hw.tag_1210.q;
  assign rcache_line[4][186].tag_reg.qe       = reg2hw.tag_1210.qe;
  assign rcache_line[4][186].tag_reg.re       = reg2hw.tag_1210.re;
  assign rcache_line[4][186].status_reg.status = reg2hw.status_1210.q;//status_reg_t'(reg2hw.status_1210.q);
  assign rcache_line[4][186].status_reg.qe    = reg2hw.status_1210.qe;
  assign rcache_line[4][186].status_reg.re    = reg2hw.status_1210.re;


  assign rcache_line[4][187].tag_reg.tag      = reg2hw.tag_1211.q;
  assign rcache_line[4][187].tag_reg.qe       = reg2hw.tag_1211.qe;
  assign rcache_line[4][187].tag_reg.re       = reg2hw.tag_1211.re;
  assign rcache_line[4][187].status_reg.status = reg2hw.status_1211.q;//status_reg_t'(reg2hw.status_1211.q);
  assign rcache_line[4][187].status_reg.qe    = reg2hw.status_1211.qe;
  assign rcache_line[4][187].status_reg.re    = reg2hw.status_1211.re;


  assign rcache_line[4][188].tag_reg.tag      = reg2hw.tag_1212.q;
  assign rcache_line[4][188].tag_reg.qe       = reg2hw.tag_1212.qe;
  assign rcache_line[4][188].tag_reg.re       = reg2hw.tag_1212.re;
  assign rcache_line[4][188].status_reg.status = reg2hw.status_1212.q;//status_reg_t'(reg2hw.status_1212.q);
  assign rcache_line[4][188].status_reg.qe    = reg2hw.status_1212.qe;
  assign rcache_line[4][188].status_reg.re    = reg2hw.status_1212.re;


  assign rcache_line[4][189].tag_reg.tag      = reg2hw.tag_1213.q;
  assign rcache_line[4][189].tag_reg.qe       = reg2hw.tag_1213.qe;
  assign rcache_line[4][189].tag_reg.re       = reg2hw.tag_1213.re;
  assign rcache_line[4][189].status_reg.status = reg2hw.status_1213.q;//status_reg_t'(reg2hw.status_1213.q);
  assign rcache_line[4][189].status_reg.qe    = reg2hw.status_1213.qe;
  assign rcache_line[4][189].status_reg.re    = reg2hw.status_1213.re;


  assign rcache_line[4][190].tag_reg.tag      = reg2hw.tag_1214.q;
  assign rcache_line[4][190].tag_reg.qe       = reg2hw.tag_1214.qe;
  assign rcache_line[4][190].tag_reg.re       = reg2hw.tag_1214.re;
  assign rcache_line[4][190].status_reg.status = reg2hw.status_1214.q;//status_reg_t'(reg2hw.status_1214.q);
  assign rcache_line[4][190].status_reg.qe    = reg2hw.status_1214.qe;
  assign rcache_line[4][190].status_reg.re    = reg2hw.status_1214.re;


  assign rcache_line[4][191].tag_reg.tag      = reg2hw.tag_1215.q;
  assign rcache_line[4][191].tag_reg.qe       = reg2hw.tag_1215.qe;
  assign rcache_line[4][191].tag_reg.re       = reg2hw.tag_1215.re;
  assign rcache_line[4][191].status_reg.status = reg2hw.status_1215.q;//status_reg_t'(reg2hw.status_1215.q);
  assign rcache_line[4][191].status_reg.qe    = reg2hw.status_1215.qe;
  assign rcache_line[4][191].status_reg.re    = reg2hw.status_1215.re;


  assign rcache_line[4][192].tag_reg.tag      = reg2hw.tag_1216.q;
  assign rcache_line[4][192].tag_reg.qe       = reg2hw.tag_1216.qe;
  assign rcache_line[4][192].tag_reg.re       = reg2hw.tag_1216.re;
  assign rcache_line[4][192].status_reg.status = reg2hw.status_1216.q;//status_reg_t'(reg2hw.status_1216.q);
  assign rcache_line[4][192].status_reg.qe    = reg2hw.status_1216.qe;
  assign rcache_line[4][192].status_reg.re    = reg2hw.status_1216.re;


  assign rcache_line[4][193].tag_reg.tag      = reg2hw.tag_1217.q;
  assign rcache_line[4][193].tag_reg.qe       = reg2hw.tag_1217.qe;
  assign rcache_line[4][193].tag_reg.re       = reg2hw.tag_1217.re;
  assign rcache_line[4][193].status_reg.status = reg2hw.status_1217.q;//status_reg_t'(reg2hw.status_1217.q);
  assign rcache_line[4][193].status_reg.qe    = reg2hw.status_1217.qe;
  assign rcache_line[4][193].status_reg.re    = reg2hw.status_1217.re;


  assign rcache_line[4][194].tag_reg.tag      = reg2hw.tag_1218.q;
  assign rcache_line[4][194].tag_reg.qe       = reg2hw.tag_1218.qe;
  assign rcache_line[4][194].tag_reg.re       = reg2hw.tag_1218.re;
  assign rcache_line[4][194].status_reg.status = reg2hw.status_1218.q;//status_reg_t'(reg2hw.status_1218.q);
  assign rcache_line[4][194].status_reg.qe    = reg2hw.status_1218.qe;
  assign rcache_line[4][194].status_reg.re    = reg2hw.status_1218.re;


  assign rcache_line[4][195].tag_reg.tag      = reg2hw.tag_1219.q;
  assign rcache_line[4][195].tag_reg.qe       = reg2hw.tag_1219.qe;
  assign rcache_line[4][195].tag_reg.re       = reg2hw.tag_1219.re;
  assign rcache_line[4][195].status_reg.status = reg2hw.status_1219.q;//status_reg_t'(reg2hw.status_1219.q);
  assign rcache_line[4][195].status_reg.qe    = reg2hw.status_1219.qe;
  assign rcache_line[4][195].status_reg.re    = reg2hw.status_1219.re;


  assign rcache_line[4][196].tag_reg.tag      = reg2hw.tag_1220.q;
  assign rcache_line[4][196].tag_reg.qe       = reg2hw.tag_1220.qe;
  assign rcache_line[4][196].tag_reg.re       = reg2hw.tag_1220.re;
  assign rcache_line[4][196].status_reg.status = reg2hw.status_1220.q;//status_reg_t'(reg2hw.status_1220.q);
  assign rcache_line[4][196].status_reg.qe    = reg2hw.status_1220.qe;
  assign rcache_line[4][196].status_reg.re    = reg2hw.status_1220.re;


  assign rcache_line[4][197].tag_reg.tag      = reg2hw.tag_1221.q;
  assign rcache_line[4][197].tag_reg.qe       = reg2hw.tag_1221.qe;
  assign rcache_line[4][197].tag_reg.re       = reg2hw.tag_1221.re;
  assign rcache_line[4][197].status_reg.status = reg2hw.status_1221.q;//status_reg_t'(reg2hw.status_1221.q);
  assign rcache_line[4][197].status_reg.qe    = reg2hw.status_1221.qe;
  assign rcache_line[4][197].status_reg.re    = reg2hw.status_1221.re;


  assign rcache_line[4][198].tag_reg.tag      = reg2hw.tag_1222.q;
  assign rcache_line[4][198].tag_reg.qe       = reg2hw.tag_1222.qe;
  assign rcache_line[4][198].tag_reg.re       = reg2hw.tag_1222.re;
  assign rcache_line[4][198].status_reg.status = reg2hw.status_1222.q;//status_reg_t'(reg2hw.status_1222.q);
  assign rcache_line[4][198].status_reg.qe    = reg2hw.status_1222.qe;
  assign rcache_line[4][198].status_reg.re    = reg2hw.status_1222.re;


  assign rcache_line[4][199].tag_reg.tag      = reg2hw.tag_1223.q;
  assign rcache_line[4][199].tag_reg.qe       = reg2hw.tag_1223.qe;
  assign rcache_line[4][199].tag_reg.re       = reg2hw.tag_1223.re;
  assign rcache_line[4][199].status_reg.status = reg2hw.status_1223.q;//status_reg_t'(reg2hw.status_1223.q);
  assign rcache_line[4][199].status_reg.qe    = reg2hw.status_1223.qe;
  assign rcache_line[4][199].status_reg.re    = reg2hw.status_1223.re;


  assign rcache_line[4][200].tag_reg.tag      = reg2hw.tag_1224.q;
  assign rcache_line[4][200].tag_reg.qe       = reg2hw.tag_1224.qe;
  assign rcache_line[4][200].tag_reg.re       = reg2hw.tag_1224.re;
  assign rcache_line[4][200].status_reg.status = reg2hw.status_1224.q;//status_reg_t'(reg2hw.status_1224.q);
  assign rcache_line[4][200].status_reg.qe    = reg2hw.status_1224.qe;
  assign rcache_line[4][200].status_reg.re    = reg2hw.status_1224.re;


  assign rcache_line[4][201].tag_reg.tag      = reg2hw.tag_1225.q;
  assign rcache_line[4][201].tag_reg.qe       = reg2hw.tag_1225.qe;
  assign rcache_line[4][201].tag_reg.re       = reg2hw.tag_1225.re;
  assign rcache_line[4][201].status_reg.status = reg2hw.status_1225.q;//status_reg_t'(reg2hw.status_1225.q);
  assign rcache_line[4][201].status_reg.qe    = reg2hw.status_1225.qe;
  assign rcache_line[4][201].status_reg.re    = reg2hw.status_1225.re;


  assign rcache_line[4][202].tag_reg.tag      = reg2hw.tag_1226.q;
  assign rcache_line[4][202].tag_reg.qe       = reg2hw.tag_1226.qe;
  assign rcache_line[4][202].tag_reg.re       = reg2hw.tag_1226.re;
  assign rcache_line[4][202].status_reg.status = reg2hw.status_1226.q;//status_reg_t'(reg2hw.status_1226.q);
  assign rcache_line[4][202].status_reg.qe    = reg2hw.status_1226.qe;
  assign rcache_line[4][202].status_reg.re    = reg2hw.status_1226.re;


  assign rcache_line[4][203].tag_reg.tag      = reg2hw.tag_1227.q;
  assign rcache_line[4][203].tag_reg.qe       = reg2hw.tag_1227.qe;
  assign rcache_line[4][203].tag_reg.re       = reg2hw.tag_1227.re;
  assign rcache_line[4][203].status_reg.status = reg2hw.status_1227.q;//status_reg_t'(reg2hw.status_1227.q);
  assign rcache_line[4][203].status_reg.qe    = reg2hw.status_1227.qe;
  assign rcache_line[4][203].status_reg.re    = reg2hw.status_1227.re;


  assign rcache_line[4][204].tag_reg.tag      = reg2hw.tag_1228.q;
  assign rcache_line[4][204].tag_reg.qe       = reg2hw.tag_1228.qe;
  assign rcache_line[4][204].tag_reg.re       = reg2hw.tag_1228.re;
  assign rcache_line[4][204].status_reg.status = reg2hw.status_1228.q;//status_reg_t'(reg2hw.status_1228.q);
  assign rcache_line[4][204].status_reg.qe    = reg2hw.status_1228.qe;
  assign rcache_line[4][204].status_reg.re    = reg2hw.status_1228.re;


  assign rcache_line[4][205].tag_reg.tag      = reg2hw.tag_1229.q;
  assign rcache_line[4][205].tag_reg.qe       = reg2hw.tag_1229.qe;
  assign rcache_line[4][205].tag_reg.re       = reg2hw.tag_1229.re;
  assign rcache_line[4][205].status_reg.status = reg2hw.status_1229.q;//status_reg_t'(reg2hw.status_1229.q);
  assign rcache_line[4][205].status_reg.qe    = reg2hw.status_1229.qe;
  assign rcache_line[4][205].status_reg.re    = reg2hw.status_1229.re;


  assign rcache_line[4][206].tag_reg.tag      = reg2hw.tag_1230.q;
  assign rcache_line[4][206].tag_reg.qe       = reg2hw.tag_1230.qe;
  assign rcache_line[4][206].tag_reg.re       = reg2hw.tag_1230.re;
  assign rcache_line[4][206].status_reg.status = reg2hw.status_1230.q;//status_reg_t'(reg2hw.status_1230.q);
  assign rcache_line[4][206].status_reg.qe    = reg2hw.status_1230.qe;
  assign rcache_line[4][206].status_reg.re    = reg2hw.status_1230.re;


  assign rcache_line[4][207].tag_reg.tag      = reg2hw.tag_1231.q;
  assign rcache_line[4][207].tag_reg.qe       = reg2hw.tag_1231.qe;
  assign rcache_line[4][207].tag_reg.re       = reg2hw.tag_1231.re;
  assign rcache_line[4][207].status_reg.status = reg2hw.status_1231.q;//status_reg_t'(reg2hw.status_1231.q);
  assign rcache_line[4][207].status_reg.qe    = reg2hw.status_1231.qe;
  assign rcache_line[4][207].status_reg.re    = reg2hw.status_1231.re;


  assign rcache_line[4][208].tag_reg.tag      = reg2hw.tag_1232.q;
  assign rcache_line[4][208].tag_reg.qe       = reg2hw.tag_1232.qe;
  assign rcache_line[4][208].tag_reg.re       = reg2hw.tag_1232.re;
  assign rcache_line[4][208].status_reg.status = reg2hw.status_1232.q;//status_reg_t'(reg2hw.status_1232.q);
  assign rcache_line[4][208].status_reg.qe    = reg2hw.status_1232.qe;
  assign rcache_line[4][208].status_reg.re    = reg2hw.status_1232.re;


  assign rcache_line[4][209].tag_reg.tag      = reg2hw.tag_1233.q;
  assign rcache_line[4][209].tag_reg.qe       = reg2hw.tag_1233.qe;
  assign rcache_line[4][209].tag_reg.re       = reg2hw.tag_1233.re;
  assign rcache_line[4][209].status_reg.status = reg2hw.status_1233.q;//status_reg_t'(reg2hw.status_1233.q);
  assign rcache_line[4][209].status_reg.qe    = reg2hw.status_1233.qe;
  assign rcache_line[4][209].status_reg.re    = reg2hw.status_1233.re;


  assign rcache_line[4][210].tag_reg.tag      = reg2hw.tag_1234.q;
  assign rcache_line[4][210].tag_reg.qe       = reg2hw.tag_1234.qe;
  assign rcache_line[4][210].tag_reg.re       = reg2hw.tag_1234.re;
  assign rcache_line[4][210].status_reg.status = reg2hw.status_1234.q;//status_reg_t'(reg2hw.status_1234.q);
  assign rcache_line[4][210].status_reg.qe    = reg2hw.status_1234.qe;
  assign rcache_line[4][210].status_reg.re    = reg2hw.status_1234.re;


  assign rcache_line[4][211].tag_reg.tag      = reg2hw.tag_1235.q;
  assign rcache_line[4][211].tag_reg.qe       = reg2hw.tag_1235.qe;
  assign rcache_line[4][211].tag_reg.re       = reg2hw.tag_1235.re;
  assign rcache_line[4][211].status_reg.status = reg2hw.status_1235.q;//status_reg_t'(reg2hw.status_1235.q);
  assign rcache_line[4][211].status_reg.qe    = reg2hw.status_1235.qe;
  assign rcache_line[4][211].status_reg.re    = reg2hw.status_1235.re;


  assign rcache_line[4][212].tag_reg.tag      = reg2hw.tag_1236.q;
  assign rcache_line[4][212].tag_reg.qe       = reg2hw.tag_1236.qe;
  assign rcache_line[4][212].tag_reg.re       = reg2hw.tag_1236.re;
  assign rcache_line[4][212].status_reg.status = reg2hw.status_1236.q;//status_reg_t'(reg2hw.status_1236.q);
  assign rcache_line[4][212].status_reg.qe    = reg2hw.status_1236.qe;
  assign rcache_line[4][212].status_reg.re    = reg2hw.status_1236.re;


  assign rcache_line[4][213].tag_reg.tag      = reg2hw.tag_1237.q;
  assign rcache_line[4][213].tag_reg.qe       = reg2hw.tag_1237.qe;
  assign rcache_line[4][213].tag_reg.re       = reg2hw.tag_1237.re;
  assign rcache_line[4][213].status_reg.status = reg2hw.status_1237.q;//status_reg_t'(reg2hw.status_1237.q);
  assign rcache_line[4][213].status_reg.qe    = reg2hw.status_1237.qe;
  assign rcache_line[4][213].status_reg.re    = reg2hw.status_1237.re;


  assign rcache_line[4][214].tag_reg.tag      = reg2hw.tag_1238.q;
  assign rcache_line[4][214].tag_reg.qe       = reg2hw.tag_1238.qe;
  assign rcache_line[4][214].tag_reg.re       = reg2hw.tag_1238.re;
  assign rcache_line[4][214].status_reg.status = reg2hw.status_1238.q;//status_reg_t'(reg2hw.status_1238.q);
  assign rcache_line[4][214].status_reg.qe    = reg2hw.status_1238.qe;
  assign rcache_line[4][214].status_reg.re    = reg2hw.status_1238.re;


  assign rcache_line[4][215].tag_reg.tag      = reg2hw.tag_1239.q;
  assign rcache_line[4][215].tag_reg.qe       = reg2hw.tag_1239.qe;
  assign rcache_line[4][215].tag_reg.re       = reg2hw.tag_1239.re;
  assign rcache_line[4][215].status_reg.status = reg2hw.status_1239.q;//status_reg_t'(reg2hw.status_1239.q);
  assign rcache_line[4][215].status_reg.qe    = reg2hw.status_1239.qe;
  assign rcache_line[4][215].status_reg.re    = reg2hw.status_1239.re;


  assign rcache_line[4][216].tag_reg.tag      = reg2hw.tag_1240.q;
  assign rcache_line[4][216].tag_reg.qe       = reg2hw.tag_1240.qe;
  assign rcache_line[4][216].tag_reg.re       = reg2hw.tag_1240.re;
  assign rcache_line[4][216].status_reg.status = reg2hw.status_1240.q;//status_reg_t'(reg2hw.status_1240.q);
  assign rcache_line[4][216].status_reg.qe    = reg2hw.status_1240.qe;
  assign rcache_line[4][216].status_reg.re    = reg2hw.status_1240.re;


  assign rcache_line[4][217].tag_reg.tag      = reg2hw.tag_1241.q;
  assign rcache_line[4][217].tag_reg.qe       = reg2hw.tag_1241.qe;
  assign rcache_line[4][217].tag_reg.re       = reg2hw.tag_1241.re;
  assign rcache_line[4][217].status_reg.status = reg2hw.status_1241.q;//status_reg_t'(reg2hw.status_1241.q);
  assign rcache_line[4][217].status_reg.qe    = reg2hw.status_1241.qe;
  assign rcache_line[4][217].status_reg.re    = reg2hw.status_1241.re;


  assign rcache_line[4][218].tag_reg.tag      = reg2hw.tag_1242.q;
  assign rcache_line[4][218].tag_reg.qe       = reg2hw.tag_1242.qe;
  assign rcache_line[4][218].tag_reg.re       = reg2hw.tag_1242.re;
  assign rcache_line[4][218].status_reg.status = reg2hw.status_1242.q;//status_reg_t'(reg2hw.status_1242.q);
  assign rcache_line[4][218].status_reg.qe    = reg2hw.status_1242.qe;
  assign rcache_line[4][218].status_reg.re    = reg2hw.status_1242.re;


  assign rcache_line[4][219].tag_reg.tag      = reg2hw.tag_1243.q;
  assign rcache_line[4][219].tag_reg.qe       = reg2hw.tag_1243.qe;
  assign rcache_line[4][219].tag_reg.re       = reg2hw.tag_1243.re;
  assign rcache_line[4][219].status_reg.status = reg2hw.status_1243.q;//status_reg_t'(reg2hw.status_1243.q);
  assign rcache_line[4][219].status_reg.qe    = reg2hw.status_1243.qe;
  assign rcache_line[4][219].status_reg.re    = reg2hw.status_1243.re;


  assign rcache_line[4][220].tag_reg.tag      = reg2hw.tag_1244.q;
  assign rcache_line[4][220].tag_reg.qe       = reg2hw.tag_1244.qe;
  assign rcache_line[4][220].tag_reg.re       = reg2hw.tag_1244.re;
  assign rcache_line[4][220].status_reg.status = reg2hw.status_1244.q;//status_reg_t'(reg2hw.status_1244.q);
  assign rcache_line[4][220].status_reg.qe    = reg2hw.status_1244.qe;
  assign rcache_line[4][220].status_reg.re    = reg2hw.status_1244.re;


  assign rcache_line[4][221].tag_reg.tag      = reg2hw.tag_1245.q;
  assign rcache_line[4][221].tag_reg.qe       = reg2hw.tag_1245.qe;
  assign rcache_line[4][221].tag_reg.re       = reg2hw.tag_1245.re;
  assign rcache_line[4][221].status_reg.status = reg2hw.status_1245.q;//status_reg_t'(reg2hw.status_1245.q);
  assign rcache_line[4][221].status_reg.qe    = reg2hw.status_1245.qe;
  assign rcache_line[4][221].status_reg.re    = reg2hw.status_1245.re;


  assign rcache_line[4][222].tag_reg.tag      = reg2hw.tag_1246.q;
  assign rcache_line[4][222].tag_reg.qe       = reg2hw.tag_1246.qe;
  assign rcache_line[4][222].tag_reg.re       = reg2hw.tag_1246.re;
  assign rcache_line[4][222].status_reg.status = reg2hw.status_1246.q;//status_reg_t'(reg2hw.status_1246.q);
  assign rcache_line[4][222].status_reg.qe    = reg2hw.status_1246.qe;
  assign rcache_line[4][222].status_reg.re    = reg2hw.status_1246.re;


  assign rcache_line[4][223].tag_reg.tag      = reg2hw.tag_1247.q;
  assign rcache_line[4][223].tag_reg.qe       = reg2hw.tag_1247.qe;
  assign rcache_line[4][223].tag_reg.re       = reg2hw.tag_1247.re;
  assign rcache_line[4][223].status_reg.status = reg2hw.status_1247.q;//status_reg_t'(reg2hw.status_1247.q);
  assign rcache_line[4][223].status_reg.qe    = reg2hw.status_1247.qe;
  assign rcache_line[4][223].status_reg.re    = reg2hw.status_1247.re;


  assign rcache_line[4][224].tag_reg.tag      = reg2hw.tag_1248.q;
  assign rcache_line[4][224].tag_reg.qe       = reg2hw.tag_1248.qe;
  assign rcache_line[4][224].tag_reg.re       = reg2hw.tag_1248.re;
  assign rcache_line[4][224].status_reg.status = reg2hw.status_1248.q;//status_reg_t'(reg2hw.status_1248.q);
  assign rcache_line[4][224].status_reg.qe    = reg2hw.status_1248.qe;
  assign rcache_line[4][224].status_reg.re    = reg2hw.status_1248.re;


  assign rcache_line[4][225].tag_reg.tag      = reg2hw.tag_1249.q;
  assign rcache_line[4][225].tag_reg.qe       = reg2hw.tag_1249.qe;
  assign rcache_line[4][225].tag_reg.re       = reg2hw.tag_1249.re;
  assign rcache_line[4][225].status_reg.status = reg2hw.status_1249.q;//status_reg_t'(reg2hw.status_1249.q);
  assign rcache_line[4][225].status_reg.qe    = reg2hw.status_1249.qe;
  assign rcache_line[4][225].status_reg.re    = reg2hw.status_1249.re;


  assign rcache_line[4][226].tag_reg.tag      = reg2hw.tag_1250.q;
  assign rcache_line[4][226].tag_reg.qe       = reg2hw.tag_1250.qe;
  assign rcache_line[4][226].tag_reg.re       = reg2hw.tag_1250.re;
  assign rcache_line[4][226].status_reg.status = reg2hw.status_1250.q;//status_reg_t'(reg2hw.status_1250.q);
  assign rcache_line[4][226].status_reg.qe    = reg2hw.status_1250.qe;
  assign rcache_line[4][226].status_reg.re    = reg2hw.status_1250.re;


  assign rcache_line[4][227].tag_reg.tag      = reg2hw.tag_1251.q;
  assign rcache_line[4][227].tag_reg.qe       = reg2hw.tag_1251.qe;
  assign rcache_line[4][227].tag_reg.re       = reg2hw.tag_1251.re;
  assign rcache_line[4][227].status_reg.status = reg2hw.status_1251.q;//status_reg_t'(reg2hw.status_1251.q);
  assign rcache_line[4][227].status_reg.qe    = reg2hw.status_1251.qe;
  assign rcache_line[4][227].status_reg.re    = reg2hw.status_1251.re;


  assign rcache_line[4][228].tag_reg.tag      = reg2hw.tag_1252.q;
  assign rcache_line[4][228].tag_reg.qe       = reg2hw.tag_1252.qe;
  assign rcache_line[4][228].tag_reg.re       = reg2hw.tag_1252.re;
  assign rcache_line[4][228].status_reg.status = reg2hw.status_1252.q;//status_reg_t'(reg2hw.status_1252.q);
  assign rcache_line[4][228].status_reg.qe    = reg2hw.status_1252.qe;
  assign rcache_line[4][228].status_reg.re    = reg2hw.status_1252.re;


  assign rcache_line[4][229].tag_reg.tag      = reg2hw.tag_1253.q;
  assign rcache_line[4][229].tag_reg.qe       = reg2hw.tag_1253.qe;
  assign rcache_line[4][229].tag_reg.re       = reg2hw.tag_1253.re;
  assign rcache_line[4][229].status_reg.status = reg2hw.status_1253.q;//status_reg_t'(reg2hw.status_1253.q);
  assign rcache_line[4][229].status_reg.qe    = reg2hw.status_1253.qe;
  assign rcache_line[4][229].status_reg.re    = reg2hw.status_1253.re;


  assign rcache_line[4][230].tag_reg.tag      = reg2hw.tag_1254.q;
  assign rcache_line[4][230].tag_reg.qe       = reg2hw.tag_1254.qe;
  assign rcache_line[4][230].tag_reg.re       = reg2hw.tag_1254.re;
  assign rcache_line[4][230].status_reg.status = reg2hw.status_1254.q;//status_reg_t'(reg2hw.status_1254.q);
  assign rcache_line[4][230].status_reg.qe    = reg2hw.status_1254.qe;
  assign rcache_line[4][230].status_reg.re    = reg2hw.status_1254.re;


  assign rcache_line[4][231].tag_reg.tag      = reg2hw.tag_1255.q;
  assign rcache_line[4][231].tag_reg.qe       = reg2hw.tag_1255.qe;
  assign rcache_line[4][231].tag_reg.re       = reg2hw.tag_1255.re;
  assign rcache_line[4][231].status_reg.status = reg2hw.status_1255.q;//status_reg_t'(reg2hw.status_1255.q);
  assign rcache_line[4][231].status_reg.qe    = reg2hw.status_1255.qe;
  assign rcache_line[4][231].status_reg.re    = reg2hw.status_1255.re;


  assign rcache_line[4][232].tag_reg.tag      = reg2hw.tag_1256.q;
  assign rcache_line[4][232].tag_reg.qe       = reg2hw.tag_1256.qe;
  assign rcache_line[4][232].tag_reg.re       = reg2hw.tag_1256.re;
  assign rcache_line[4][232].status_reg.status = reg2hw.status_1256.q;//status_reg_t'(reg2hw.status_1256.q);
  assign rcache_line[4][232].status_reg.qe    = reg2hw.status_1256.qe;
  assign rcache_line[4][232].status_reg.re    = reg2hw.status_1256.re;


  assign rcache_line[4][233].tag_reg.tag      = reg2hw.tag_1257.q;
  assign rcache_line[4][233].tag_reg.qe       = reg2hw.tag_1257.qe;
  assign rcache_line[4][233].tag_reg.re       = reg2hw.tag_1257.re;
  assign rcache_line[4][233].status_reg.status = reg2hw.status_1257.q;//status_reg_t'(reg2hw.status_1257.q);
  assign rcache_line[4][233].status_reg.qe    = reg2hw.status_1257.qe;
  assign rcache_line[4][233].status_reg.re    = reg2hw.status_1257.re;


  assign rcache_line[4][234].tag_reg.tag      = reg2hw.tag_1258.q;
  assign rcache_line[4][234].tag_reg.qe       = reg2hw.tag_1258.qe;
  assign rcache_line[4][234].tag_reg.re       = reg2hw.tag_1258.re;
  assign rcache_line[4][234].status_reg.status = reg2hw.status_1258.q;//status_reg_t'(reg2hw.status_1258.q);
  assign rcache_line[4][234].status_reg.qe    = reg2hw.status_1258.qe;
  assign rcache_line[4][234].status_reg.re    = reg2hw.status_1258.re;


  assign rcache_line[4][235].tag_reg.tag      = reg2hw.tag_1259.q;
  assign rcache_line[4][235].tag_reg.qe       = reg2hw.tag_1259.qe;
  assign rcache_line[4][235].tag_reg.re       = reg2hw.tag_1259.re;
  assign rcache_line[4][235].status_reg.status = reg2hw.status_1259.q;//status_reg_t'(reg2hw.status_1259.q);
  assign rcache_line[4][235].status_reg.qe    = reg2hw.status_1259.qe;
  assign rcache_line[4][235].status_reg.re    = reg2hw.status_1259.re;


  assign rcache_line[4][236].tag_reg.tag      = reg2hw.tag_1260.q;
  assign rcache_line[4][236].tag_reg.qe       = reg2hw.tag_1260.qe;
  assign rcache_line[4][236].tag_reg.re       = reg2hw.tag_1260.re;
  assign rcache_line[4][236].status_reg.status = reg2hw.status_1260.q;//status_reg_t'(reg2hw.status_1260.q);
  assign rcache_line[4][236].status_reg.qe    = reg2hw.status_1260.qe;
  assign rcache_line[4][236].status_reg.re    = reg2hw.status_1260.re;


  assign rcache_line[4][237].tag_reg.tag      = reg2hw.tag_1261.q;
  assign rcache_line[4][237].tag_reg.qe       = reg2hw.tag_1261.qe;
  assign rcache_line[4][237].tag_reg.re       = reg2hw.tag_1261.re;
  assign rcache_line[4][237].status_reg.status = reg2hw.status_1261.q;//status_reg_t'(reg2hw.status_1261.q);
  assign rcache_line[4][237].status_reg.qe    = reg2hw.status_1261.qe;
  assign rcache_line[4][237].status_reg.re    = reg2hw.status_1261.re;


  assign rcache_line[4][238].tag_reg.tag      = reg2hw.tag_1262.q;
  assign rcache_line[4][238].tag_reg.qe       = reg2hw.tag_1262.qe;
  assign rcache_line[4][238].tag_reg.re       = reg2hw.tag_1262.re;
  assign rcache_line[4][238].status_reg.status = reg2hw.status_1262.q;//status_reg_t'(reg2hw.status_1262.q);
  assign rcache_line[4][238].status_reg.qe    = reg2hw.status_1262.qe;
  assign rcache_line[4][238].status_reg.re    = reg2hw.status_1262.re;


  assign rcache_line[4][239].tag_reg.tag      = reg2hw.tag_1263.q;
  assign rcache_line[4][239].tag_reg.qe       = reg2hw.tag_1263.qe;
  assign rcache_line[4][239].tag_reg.re       = reg2hw.tag_1263.re;
  assign rcache_line[4][239].status_reg.status = reg2hw.status_1263.q;//status_reg_t'(reg2hw.status_1263.q);
  assign rcache_line[4][239].status_reg.qe    = reg2hw.status_1263.qe;
  assign rcache_line[4][239].status_reg.re    = reg2hw.status_1263.re;


  assign rcache_line[4][240].tag_reg.tag      = reg2hw.tag_1264.q;
  assign rcache_line[4][240].tag_reg.qe       = reg2hw.tag_1264.qe;
  assign rcache_line[4][240].tag_reg.re       = reg2hw.tag_1264.re;
  assign rcache_line[4][240].status_reg.status = reg2hw.status_1264.q;//status_reg_t'(reg2hw.status_1264.q);
  assign rcache_line[4][240].status_reg.qe    = reg2hw.status_1264.qe;
  assign rcache_line[4][240].status_reg.re    = reg2hw.status_1264.re;


  assign rcache_line[4][241].tag_reg.tag      = reg2hw.tag_1265.q;
  assign rcache_line[4][241].tag_reg.qe       = reg2hw.tag_1265.qe;
  assign rcache_line[4][241].tag_reg.re       = reg2hw.tag_1265.re;
  assign rcache_line[4][241].status_reg.status = reg2hw.status_1265.q;//status_reg_t'(reg2hw.status_1265.q);
  assign rcache_line[4][241].status_reg.qe    = reg2hw.status_1265.qe;
  assign rcache_line[4][241].status_reg.re    = reg2hw.status_1265.re;


  assign rcache_line[4][242].tag_reg.tag      = reg2hw.tag_1266.q;
  assign rcache_line[4][242].tag_reg.qe       = reg2hw.tag_1266.qe;
  assign rcache_line[4][242].tag_reg.re       = reg2hw.tag_1266.re;
  assign rcache_line[4][242].status_reg.status = reg2hw.status_1266.q;//status_reg_t'(reg2hw.status_1266.q);
  assign rcache_line[4][242].status_reg.qe    = reg2hw.status_1266.qe;
  assign rcache_line[4][242].status_reg.re    = reg2hw.status_1266.re;


  assign rcache_line[4][243].tag_reg.tag      = reg2hw.tag_1267.q;
  assign rcache_line[4][243].tag_reg.qe       = reg2hw.tag_1267.qe;
  assign rcache_line[4][243].tag_reg.re       = reg2hw.tag_1267.re;
  assign rcache_line[4][243].status_reg.status = reg2hw.status_1267.q;//status_reg_t'(reg2hw.status_1267.q);
  assign rcache_line[4][243].status_reg.qe    = reg2hw.status_1267.qe;
  assign rcache_line[4][243].status_reg.re    = reg2hw.status_1267.re;


  assign rcache_line[4][244].tag_reg.tag      = reg2hw.tag_1268.q;
  assign rcache_line[4][244].tag_reg.qe       = reg2hw.tag_1268.qe;
  assign rcache_line[4][244].tag_reg.re       = reg2hw.tag_1268.re;
  assign rcache_line[4][244].status_reg.status = reg2hw.status_1268.q;//status_reg_t'(reg2hw.status_1268.q);
  assign rcache_line[4][244].status_reg.qe    = reg2hw.status_1268.qe;
  assign rcache_line[4][244].status_reg.re    = reg2hw.status_1268.re;


  assign rcache_line[4][245].tag_reg.tag      = reg2hw.tag_1269.q;
  assign rcache_line[4][245].tag_reg.qe       = reg2hw.tag_1269.qe;
  assign rcache_line[4][245].tag_reg.re       = reg2hw.tag_1269.re;
  assign rcache_line[4][245].status_reg.status = reg2hw.status_1269.q;//status_reg_t'(reg2hw.status_1269.q);
  assign rcache_line[4][245].status_reg.qe    = reg2hw.status_1269.qe;
  assign rcache_line[4][245].status_reg.re    = reg2hw.status_1269.re;


  assign rcache_line[4][246].tag_reg.tag      = reg2hw.tag_1270.q;
  assign rcache_line[4][246].tag_reg.qe       = reg2hw.tag_1270.qe;
  assign rcache_line[4][246].tag_reg.re       = reg2hw.tag_1270.re;
  assign rcache_line[4][246].status_reg.status = reg2hw.status_1270.q;//status_reg_t'(reg2hw.status_1270.q);
  assign rcache_line[4][246].status_reg.qe    = reg2hw.status_1270.qe;
  assign rcache_line[4][246].status_reg.re    = reg2hw.status_1270.re;


  assign rcache_line[4][247].tag_reg.tag      = reg2hw.tag_1271.q;
  assign rcache_line[4][247].tag_reg.qe       = reg2hw.tag_1271.qe;
  assign rcache_line[4][247].tag_reg.re       = reg2hw.tag_1271.re;
  assign rcache_line[4][247].status_reg.status = reg2hw.status_1271.q;//status_reg_t'(reg2hw.status_1271.q);
  assign rcache_line[4][247].status_reg.qe    = reg2hw.status_1271.qe;
  assign rcache_line[4][247].status_reg.re    = reg2hw.status_1271.re;


  assign rcache_line[4][248].tag_reg.tag      = reg2hw.tag_1272.q;
  assign rcache_line[4][248].tag_reg.qe       = reg2hw.tag_1272.qe;
  assign rcache_line[4][248].tag_reg.re       = reg2hw.tag_1272.re;
  assign rcache_line[4][248].status_reg.status = reg2hw.status_1272.q;//status_reg_t'(reg2hw.status_1272.q);
  assign rcache_line[4][248].status_reg.qe    = reg2hw.status_1272.qe;
  assign rcache_line[4][248].status_reg.re    = reg2hw.status_1272.re;


  assign rcache_line[4][249].tag_reg.tag      = reg2hw.tag_1273.q;
  assign rcache_line[4][249].tag_reg.qe       = reg2hw.tag_1273.qe;
  assign rcache_line[4][249].tag_reg.re       = reg2hw.tag_1273.re;
  assign rcache_line[4][249].status_reg.status = reg2hw.status_1273.q;//status_reg_t'(reg2hw.status_1273.q);
  assign rcache_line[4][249].status_reg.qe    = reg2hw.status_1273.qe;
  assign rcache_line[4][249].status_reg.re    = reg2hw.status_1273.re;


  assign rcache_line[4][250].tag_reg.tag      = reg2hw.tag_1274.q;
  assign rcache_line[4][250].tag_reg.qe       = reg2hw.tag_1274.qe;
  assign rcache_line[4][250].tag_reg.re       = reg2hw.tag_1274.re;
  assign rcache_line[4][250].status_reg.status = reg2hw.status_1274.q;//status_reg_t'(reg2hw.status_1274.q);
  assign rcache_line[4][250].status_reg.qe    = reg2hw.status_1274.qe;
  assign rcache_line[4][250].status_reg.re    = reg2hw.status_1274.re;


  assign rcache_line[4][251].tag_reg.tag      = reg2hw.tag_1275.q;
  assign rcache_line[4][251].tag_reg.qe       = reg2hw.tag_1275.qe;
  assign rcache_line[4][251].tag_reg.re       = reg2hw.tag_1275.re;
  assign rcache_line[4][251].status_reg.status = reg2hw.status_1275.q;//status_reg_t'(reg2hw.status_1275.q);
  assign rcache_line[4][251].status_reg.qe    = reg2hw.status_1275.qe;
  assign rcache_line[4][251].status_reg.re    = reg2hw.status_1275.re;


  assign rcache_line[4][252].tag_reg.tag      = reg2hw.tag_1276.q;
  assign rcache_line[4][252].tag_reg.qe       = reg2hw.tag_1276.qe;
  assign rcache_line[4][252].tag_reg.re       = reg2hw.tag_1276.re;
  assign rcache_line[4][252].status_reg.status = reg2hw.status_1276.q;//status_reg_t'(reg2hw.status_1276.q);
  assign rcache_line[4][252].status_reg.qe    = reg2hw.status_1276.qe;
  assign rcache_line[4][252].status_reg.re    = reg2hw.status_1276.re;


  assign rcache_line[4][253].tag_reg.tag      = reg2hw.tag_1277.q;
  assign rcache_line[4][253].tag_reg.qe       = reg2hw.tag_1277.qe;
  assign rcache_line[4][253].tag_reg.re       = reg2hw.tag_1277.re;
  assign rcache_line[4][253].status_reg.status = reg2hw.status_1277.q;//status_reg_t'(reg2hw.status_1277.q);
  assign rcache_line[4][253].status_reg.qe    = reg2hw.status_1277.qe;
  assign rcache_line[4][253].status_reg.re    = reg2hw.status_1277.re;


  assign rcache_line[4][254].tag_reg.tag      = reg2hw.tag_1278.q;
  assign rcache_line[4][254].tag_reg.qe       = reg2hw.tag_1278.qe;
  assign rcache_line[4][254].tag_reg.re       = reg2hw.tag_1278.re;
  assign rcache_line[4][254].status_reg.status = reg2hw.status_1278.q;//status_reg_t'(reg2hw.status_1278.q);
  assign rcache_line[4][254].status_reg.qe    = reg2hw.status_1278.qe;
  assign rcache_line[4][254].status_reg.re    = reg2hw.status_1278.re;


  assign rcache_line[4][255].tag_reg.tag      = reg2hw.tag_1279.q;
  assign rcache_line[4][255].tag_reg.qe       = reg2hw.tag_1279.qe;
  assign rcache_line[4][255].tag_reg.re       = reg2hw.tag_1279.re;
  assign rcache_line[4][255].status_reg.status = reg2hw.status_1279.q;//status_reg_t'(reg2hw.status_1279.q);
  assign rcache_line[4][255].status_reg.qe    = reg2hw.status_1279.qe;
  assign rcache_line[4][255].status_reg.re    = reg2hw.status_1279.re;


  assign rcache_line[5][0].tag_reg.tag      = reg2hw.tag_1280.q;
  assign rcache_line[5][0].tag_reg.qe       = reg2hw.tag_1280.qe;
  assign rcache_line[5][0].tag_reg.re       = reg2hw.tag_1280.re;
  assign rcache_line[5][0].status_reg.status = reg2hw.status_1280.q;//status_reg_t'(reg2hw.status_1280.q);
  assign rcache_line[5][0].status_reg.qe    = reg2hw.status_1280.qe;
  assign rcache_line[5][0].status_reg.re    = reg2hw.status_1280.re;


  assign rcache_line[5][1].tag_reg.tag      = reg2hw.tag_1281.q;
  assign rcache_line[5][1].tag_reg.qe       = reg2hw.tag_1281.qe;
  assign rcache_line[5][1].tag_reg.re       = reg2hw.tag_1281.re;
  assign rcache_line[5][1].status_reg.status = reg2hw.status_1281.q;//status_reg_t'(reg2hw.status_1281.q);
  assign rcache_line[5][1].status_reg.qe    = reg2hw.status_1281.qe;
  assign rcache_line[5][1].status_reg.re    = reg2hw.status_1281.re;


  assign rcache_line[5][2].tag_reg.tag      = reg2hw.tag_1282.q;
  assign rcache_line[5][2].tag_reg.qe       = reg2hw.tag_1282.qe;
  assign rcache_line[5][2].tag_reg.re       = reg2hw.tag_1282.re;
  assign rcache_line[5][2].status_reg.status = reg2hw.status_1282.q;//status_reg_t'(reg2hw.status_1282.q);
  assign rcache_line[5][2].status_reg.qe    = reg2hw.status_1282.qe;
  assign rcache_line[5][2].status_reg.re    = reg2hw.status_1282.re;


  assign rcache_line[5][3].tag_reg.tag      = reg2hw.tag_1283.q;
  assign rcache_line[5][3].tag_reg.qe       = reg2hw.tag_1283.qe;
  assign rcache_line[5][3].tag_reg.re       = reg2hw.tag_1283.re;
  assign rcache_line[5][3].status_reg.status = reg2hw.status_1283.q;//status_reg_t'(reg2hw.status_1283.q);
  assign rcache_line[5][3].status_reg.qe    = reg2hw.status_1283.qe;
  assign rcache_line[5][3].status_reg.re    = reg2hw.status_1283.re;


  assign rcache_line[5][4].tag_reg.tag      = reg2hw.tag_1284.q;
  assign rcache_line[5][4].tag_reg.qe       = reg2hw.tag_1284.qe;
  assign rcache_line[5][4].tag_reg.re       = reg2hw.tag_1284.re;
  assign rcache_line[5][4].status_reg.status = reg2hw.status_1284.q;//status_reg_t'(reg2hw.status_1284.q);
  assign rcache_line[5][4].status_reg.qe    = reg2hw.status_1284.qe;
  assign rcache_line[5][4].status_reg.re    = reg2hw.status_1284.re;


  assign rcache_line[5][5].tag_reg.tag      = reg2hw.tag_1285.q;
  assign rcache_line[5][5].tag_reg.qe       = reg2hw.tag_1285.qe;
  assign rcache_line[5][5].tag_reg.re       = reg2hw.tag_1285.re;
  assign rcache_line[5][5].status_reg.status = reg2hw.status_1285.q;//status_reg_t'(reg2hw.status_1285.q);
  assign rcache_line[5][5].status_reg.qe    = reg2hw.status_1285.qe;
  assign rcache_line[5][5].status_reg.re    = reg2hw.status_1285.re;


  assign rcache_line[5][6].tag_reg.tag      = reg2hw.tag_1286.q;
  assign rcache_line[5][6].tag_reg.qe       = reg2hw.tag_1286.qe;
  assign rcache_line[5][6].tag_reg.re       = reg2hw.tag_1286.re;
  assign rcache_line[5][6].status_reg.status = reg2hw.status_1286.q;//status_reg_t'(reg2hw.status_1286.q);
  assign rcache_line[5][6].status_reg.qe    = reg2hw.status_1286.qe;
  assign rcache_line[5][6].status_reg.re    = reg2hw.status_1286.re;


  assign rcache_line[5][7].tag_reg.tag      = reg2hw.tag_1287.q;
  assign rcache_line[5][7].tag_reg.qe       = reg2hw.tag_1287.qe;
  assign rcache_line[5][7].tag_reg.re       = reg2hw.tag_1287.re;
  assign rcache_line[5][7].status_reg.status = reg2hw.status_1287.q;//status_reg_t'(reg2hw.status_1287.q);
  assign rcache_line[5][7].status_reg.qe    = reg2hw.status_1287.qe;
  assign rcache_line[5][7].status_reg.re    = reg2hw.status_1287.re;


  assign rcache_line[5][8].tag_reg.tag      = reg2hw.tag_1288.q;
  assign rcache_line[5][8].tag_reg.qe       = reg2hw.tag_1288.qe;
  assign rcache_line[5][8].tag_reg.re       = reg2hw.tag_1288.re;
  assign rcache_line[5][8].status_reg.status = reg2hw.status_1288.q;//status_reg_t'(reg2hw.status_1288.q);
  assign rcache_line[5][8].status_reg.qe    = reg2hw.status_1288.qe;
  assign rcache_line[5][8].status_reg.re    = reg2hw.status_1288.re;


  assign rcache_line[5][9].tag_reg.tag      = reg2hw.tag_1289.q;
  assign rcache_line[5][9].tag_reg.qe       = reg2hw.tag_1289.qe;
  assign rcache_line[5][9].tag_reg.re       = reg2hw.tag_1289.re;
  assign rcache_line[5][9].status_reg.status = reg2hw.status_1289.q;//status_reg_t'(reg2hw.status_1289.q);
  assign rcache_line[5][9].status_reg.qe    = reg2hw.status_1289.qe;
  assign rcache_line[5][9].status_reg.re    = reg2hw.status_1289.re;


  assign rcache_line[5][10].tag_reg.tag      = reg2hw.tag_1290.q;
  assign rcache_line[5][10].tag_reg.qe       = reg2hw.tag_1290.qe;
  assign rcache_line[5][10].tag_reg.re       = reg2hw.tag_1290.re;
  assign rcache_line[5][10].status_reg.status = reg2hw.status_1290.q;//status_reg_t'(reg2hw.status_1290.q);
  assign rcache_line[5][10].status_reg.qe    = reg2hw.status_1290.qe;
  assign rcache_line[5][10].status_reg.re    = reg2hw.status_1290.re;


  assign rcache_line[5][11].tag_reg.tag      = reg2hw.tag_1291.q;
  assign rcache_line[5][11].tag_reg.qe       = reg2hw.tag_1291.qe;
  assign rcache_line[5][11].tag_reg.re       = reg2hw.tag_1291.re;
  assign rcache_line[5][11].status_reg.status = reg2hw.status_1291.q;//status_reg_t'(reg2hw.status_1291.q);
  assign rcache_line[5][11].status_reg.qe    = reg2hw.status_1291.qe;
  assign rcache_line[5][11].status_reg.re    = reg2hw.status_1291.re;


  assign rcache_line[5][12].tag_reg.tag      = reg2hw.tag_1292.q;
  assign rcache_line[5][12].tag_reg.qe       = reg2hw.tag_1292.qe;
  assign rcache_line[5][12].tag_reg.re       = reg2hw.tag_1292.re;
  assign rcache_line[5][12].status_reg.status = reg2hw.status_1292.q;//status_reg_t'(reg2hw.status_1292.q);
  assign rcache_line[5][12].status_reg.qe    = reg2hw.status_1292.qe;
  assign rcache_line[5][12].status_reg.re    = reg2hw.status_1292.re;


  assign rcache_line[5][13].tag_reg.tag      = reg2hw.tag_1293.q;
  assign rcache_line[5][13].tag_reg.qe       = reg2hw.tag_1293.qe;
  assign rcache_line[5][13].tag_reg.re       = reg2hw.tag_1293.re;
  assign rcache_line[5][13].status_reg.status = reg2hw.status_1293.q;//status_reg_t'(reg2hw.status_1293.q);
  assign rcache_line[5][13].status_reg.qe    = reg2hw.status_1293.qe;
  assign rcache_line[5][13].status_reg.re    = reg2hw.status_1293.re;


  assign rcache_line[5][14].tag_reg.tag      = reg2hw.tag_1294.q;
  assign rcache_line[5][14].tag_reg.qe       = reg2hw.tag_1294.qe;
  assign rcache_line[5][14].tag_reg.re       = reg2hw.tag_1294.re;
  assign rcache_line[5][14].status_reg.status = reg2hw.status_1294.q;//status_reg_t'(reg2hw.status_1294.q);
  assign rcache_line[5][14].status_reg.qe    = reg2hw.status_1294.qe;
  assign rcache_line[5][14].status_reg.re    = reg2hw.status_1294.re;


  assign rcache_line[5][15].tag_reg.tag      = reg2hw.tag_1295.q;
  assign rcache_line[5][15].tag_reg.qe       = reg2hw.tag_1295.qe;
  assign rcache_line[5][15].tag_reg.re       = reg2hw.tag_1295.re;
  assign rcache_line[5][15].status_reg.status = reg2hw.status_1295.q;//status_reg_t'(reg2hw.status_1295.q);
  assign rcache_line[5][15].status_reg.qe    = reg2hw.status_1295.qe;
  assign rcache_line[5][15].status_reg.re    = reg2hw.status_1295.re;


  assign rcache_line[5][16].tag_reg.tag      = reg2hw.tag_1296.q;
  assign rcache_line[5][16].tag_reg.qe       = reg2hw.tag_1296.qe;
  assign rcache_line[5][16].tag_reg.re       = reg2hw.tag_1296.re;
  assign rcache_line[5][16].status_reg.status = reg2hw.status_1296.q;//status_reg_t'(reg2hw.status_1296.q);
  assign rcache_line[5][16].status_reg.qe    = reg2hw.status_1296.qe;
  assign rcache_line[5][16].status_reg.re    = reg2hw.status_1296.re;


  assign rcache_line[5][17].tag_reg.tag      = reg2hw.tag_1297.q;
  assign rcache_line[5][17].tag_reg.qe       = reg2hw.tag_1297.qe;
  assign rcache_line[5][17].tag_reg.re       = reg2hw.tag_1297.re;
  assign rcache_line[5][17].status_reg.status = reg2hw.status_1297.q;//status_reg_t'(reg2hw.status_1297.q);
  assign rcache_line[5][17].status_reg.qe    = reg2hw.status_1297.qe;
  assign rcache_line[5][17].status_reg.re    = reg2hw.status_1297.re;


  assign rcache_line[5][18].tag_reg.tag      = reg2hw.tag_1298.q;
  assign rcache_line[5][18].tag_reg.qe       = reg2hw.tag_1298.qe;
  assign rcache_line[5][18].tag_reg.re       = reg2hw.tag_1298.re;
  assign rcache_line[5][18].status_reg.status = reg2hw.status_1298.q;//status_reg_t'(reg2hw.status_1298.q);
  assign rcache_line[5][18].status_reg.qe    = reg2hw.status_1298.qe;
  assign rcache_line[5][18].status_reg.re    = reg2hw.status_1298.re;


  assign rcache_line[5][19].tag_reg.tag      = reg2hw.tag_1299.q;
  assign rcache_line[5][19].tag_reg.qe       = reg2hw.tag_1299.qe;
  assign rcache_line[5][19].tag_reg.re       = reg2hw.tag_1299.re;
  assign rcache_line[5][19].status_reg.status = reg2hw.status_1299.q;//status_reg_t'(reg2hw.status_1299.q);
  assign rcache_line[5][19].status_reg.qe    = reg2hw.status_1299.qe;
  assign rcache_line[5][19].status_reg.re    = reg2hw.status_1299.re;


  assign rcache_line[5][20].tag_reg.tag      = reg2hw.tag_1300.q;
  assign rcache_line[5][20].tag_reg.qe       = reg2hw.tag_1300.qe;
  assign rcache_line[5][20].tag_reg.re       = reg2hw.tag_1300.re;
  assign rcache_line[5][20].status_reg.status = reg2hw.status_1300.q;//status_reg_t'(reg2hw.status_1300.q);
  assign rcache_line[5][20].status_reg.qe    = reg2hw.status_1300.qe;
  assign rcache_line[5][20].status_reg.re    = reg2hw.status_1300.re;


  assign rcache_line[5][21].tag_reg.tag      = reg2hw.tag_1301.q;
  assign rcache_line[5][21].tag_reg.qe       = reg2hw.tag_1301.qe;
  assign rcache_line[5][21].tag_reg.re       = reg2hw.tag_1301.re;
  assign rcache_line[5][21].status_reg.status = reg2hw.status_1301.q;//status_reg_t'(reg2hw.status_1301.q);
  assign rcache_line[5][21].status_reg.qe    = reg2hw.status_1301.qe;
  assign rcache_line[5][21].status_reg.re    = reg2hw.status_1301.re;


  assign rcache_line[5][22].tag_reg.tag      = reg2hw.tag_1302.q;
  assign rcache_line[5][22].tag_reg.qe       = reg2hw.tag_1302.qe;
  assign rcache_line[5][22].tag_reg.re       = reg2hw.tag_1302.re;
  assign rcache_line[5][22].status_reg.status = reg2hw.status_1302.q;//status_reg_t'(reg2hw.status_1302.q);
  assign rcache_line[5][22].status_reg.qe    = reg2hw.status_1302.qe;
  assign rcache_line[5][22].status_reg.re    = reg2hw.status_1302.re;


  assign rcache_line[5][23].tag_reg.tag      = reg2hw.tag_1303.q;
  assign rcache_line[5][23].tag_reg.qe       = reg2hw.tag_1303.qe;
  assign rcache_line[5][23].tag_reg.re       = reg2hw.tag_1303.re;
  assign rcache_line[5][23].status_reg.status = reg2hw.status_1303.q;//status_reg_t'(reg2hw.status_1303.q);
  assign rcache_line[5][23].status_reg.qe    = reg2hw.status_1303.qe;
  assign rcache_line[5][23].status_reg.re    = reg2hw.status_1303.re;


  assign rcache_line[5][24].tag_reg.tag      = reg2hw.tag_1304.q;
  assign rcache_line[5][24].tag_reg.qe       = reg2hw.tag_1304.qe;
  assign rcache_line[5][24].tag_reg.re       = reg2hw.tag_1304.re;
  assign rcache_line[5][24].status_reg.status = reg2hw.status_1304.q;//status_reg_t'(reg2hw.status_1304.q);
  assign rcache_line[5][24].status_reg.qe    = reg2hw.status_1304.qe;
  assign rcache_line[5][24].status_reg.re    = reg2hw.status_1304.re;


  assign rcache_line[5][25].tag_reg.tag      = reg2hw.tag_1305.q;
  assign rcache_line[5][25].tag_reg.qe       = reg2hw.tag_1305.qe;
  assign rcache_line[5][25].tag_reg.re       = reg2hw.tag_1305.re;
  assign rcache_line[5][25].status_reg.status = reg2hw.status_1305.q;//status_reg_t'(reg2hw.status_1305.q);
  assign rcache_line[5][25].status_reg.qe    = reg2hw.status_1305.qe;
  assign rcache_line[5][25].status_reg.re    = reg2hw.status_1305.re;


  assign rcache_line[5][26].tag_reg.tag      = reg2hw.tag_1306.q;
  assign rcache_line[5][26].tag_reg.qe       = reg2hw.tag_1306.qe;
  assign rcache_line[5][26].tag_reg.re       = reg2hw.tag_1306.re;
  assign rcache_line[5][26].status_reg.status = reg2hw.status_1306.q;//status_reg_t'(reg2hw.status_1306.q);
  assign rcache_line[5][26].status_reg.qe    = reg2hw.status_1306.qe;
  assign rcache_line[5][26].status_reg.re    = reg2hw.status_1306.re;


  assign rcache_line[5][27].tag_reg.tag      = reg2hw.tag_1307.q;
  assign rcache_line[5][27].tag_reg.qe       = reg2hw.tag_1307.qe;
  assign rcache_line[5][27].tag_reg.re       = reg2hw.tag_1307.re;
  assign rcache_line[5][27].status_reg.status = reg2hw.status_1307.q;//status_reg_t'(reg2hw.status_1307.q);
  assign rcache_line[5][27].status_reg.qe    = reg2hw.status_1307.qe;
  assign rcache_line[5][27].status_reg.re    = reg2hw.status_1307.re;


  assign rcache_line[5][28].tag_reg.tag      = reg2hw.tag_1308.q;
  assign rcache_line[5][28].tag_reg.qe       = reg2hw.tag_1308.qe;
  assign rcache_line[5][28].tag_reg.re       = reg2hw.tag_1308.re;
  assign rcache_line[5][28].status_reg.status = reg2hw.status_1308.q;//status_reg_t'(reg2hw.status_1308.q);
  assign rcache_line[5][28].status_reg.qe    = reg2hw.status_1308.qe;
  assign rcache_line[5][28].status_reg.re    = reg2hw.status_1308.re;


  assign rcache_line[5][29].tag_reg.tag      = reg2hw.tag_1309.q;
  assign rcache_line[5][29].tag_reg.qe       = reg2hw.tag_1309.qe;
  assign rcache_line[5][29].tag_reg.re       = reg2hw.tag_1309.re;
  assign rcache_line[5][29].status_reg.status = reg2hw.status_1309.q;//status_reg_t'(reg2hw.status_1309.q);
  assign rcache_line[5][29].status_reg.qe    = reg2hw.status_1309.qe;
  assign rcache_line[5][29].status_reg.re    = reg2hw.status_1309.re;


  assign rcache_line[5][30].tag_reg.tag      = reg2hw.tag_1310.q;
  assign rcache_line[5][30].tag_reg.qe       = reg2hw.tag_1310.qe;
  assign rcache_line[5][30].tag_reg.re       = reg2hw.tag_1310.re;
  assign rcache_line[5][30].status_reg.status = reg2hw.status_1310.q;//status_reg_t'(reg2hw.status_1310.q);
  assign rcache_line[5][30].status_reg.qe    = reg2hw.status_1310.qe;
  assign rcache_line[5][30].status_reg.re    = reg2hw.status_1310.re;


  assign rcache_line[5][31].tag_reg.tag      = reg2hw.tag_1311.q;
  assign rcache_line[5][31].tag_reg.qe       = reg2hw.tag_1311.qe;
  assign rcache_line[5][31].tag_reg.re       = reg2hw.tag_1311.re;
  assign rcache_line[5][31].status_reg.status = reg2hw.status_1311.q;//status_reg_t'(reg2hw.status_1311.q);
  assign rcache_line[5][31].status_reg.qe    = reg2hw.status_1311.qe;
  assign rcache_line[5][31].status_reg.re    = reg2hw.status_1311.re;


  assign rcache_line[5][32].tag_reg.tag      = reg2hw.tag_1312.q;
  assign rcache_line[5][32].tag_reg.qe       = reg2hw.tag_1312.qe;
  assign rcache_line[5][32].tag_reg.re       = reg2hw.tag_1312.re;
  assign rcache_line[5][32].status_reg.status = reg2hw.status_1312.q;//status_reg_t'(reg2hw.status_1312.q);
  assign rcache_line[5][32].status_reg.qe    = reg2hw.status_1312.qe;
  assign rcache_line[5][32].status_reg.re    = reg2hw.status_1312.re;


  assign rcache_line[5][33].tag_reg.tag      = reg2hw.tag_1313.q;
  assign rcache_line[5][33].tag_reg.qe       = reg2hw.tag_1313.qe;
  assign rcache_line[5][33].tag_reg.re       = reg2hw.tag_1313.re;
  assign rcache_line[5][33].status_reg.status = reg2hw.status_1313.q;//status_reg_t'(reg2hw.status_1313.q);
  assign rcache_line[5][33].status_reg.qe    = reg2hw.status_1313.qe;
  assign rcache_line[5][33].status_reg.re    = reg2hw.status_1313.re;


  assign rcache_line[5][34].tag_reg.tag      = reg2hw.tag_1314.q;
  assign rcache_line[5][34].tag_reg.qe       = reg2hw.tag_1314.qe;
  assign rcache_line[5][34].tag_reg.re       = reg2hw.tag_1314.re;
  assign rcache_line[5][34].status_reg.status = reg2hw.status_1314.q;//status_reg_t'(reg2hw.status_1314.q);
  assign rcache_line[5][34].status_reg.qe    = reg2hw.status_1314.qe;
  assign rcache_line[5][34].status_reg.re    = reg2hw.status_1314.re;


  assign rcache_line[5][35].tag_reg.tag      = reg2hw.tag_1315.q;
  assign rcache_line[5][35].tag_reg.qe       = reg2hw.tag_1315.qe;
  assign rcache_line[5][35].tag_reg.re       = reg2hw.tag_1315.re;
  assign rcache_line[5][35].status_reg.status = reg2hw.status_1315.q;//status_reg_t'(reg2hw.status_1315.q);
  assign rcache_line[5][35].status_reg.qe    = reg2hw.status_1315.qe;
  assign rcache_line[5][35].status_reg.re    = reg2hw.status_1315.re;


  assign rcache_line[5][36].tag_reg.tag      = reg2hw.tag_1316.q;
  assign rcache_line[5][36].tag_reg.qe       = reg2hw.tag_1316.qe;
  assign rcache_line[5][36].tag_reg.re       = reg2hw.tag_1316.re;
  assign rcache_line[5][36].status_reg.status = reg2hw.status_1316.q;//status_reg_t'(reg2hw.status_1316.q);
  assign rcache_line[5][36].status_reg.qe    = reg2hw.status_1316.qe;
  assign rcache_line[5][36].status_reg.re    = reg2hw.status_1316.re;


  assign rcache_line[5][37].tag_reg.tag      = reg2hw.tag_1317.q;
  assign rcache_line[5][37].tag_reg.qe       = reg2hw.tag_1317.qe;
  assign rcache_line[5][37].tag_reg.re       = reg2hw.tag_1317.re;
  assign rcache_line[5][37].status_reg.status = reg2hw.status_1317.q;//status_reg_t'(reg2hw.status_1317.q);
  assign rcache_line[5][37].status_reg.qe    = reg2hw.status_1317.qe;
  assign rcache_line[5][37].status_reg.re    = reg2hw.status_1317.re;


  assign rcache_line[5][38].tag_reg.tag      = reg2hw.tag_1318.q;
  assign rcache_line[5][38].tag_reg.qe       = reg2hw.tag_1318.qe;
  assign rcache_line[5][38].tag_reg.re       = reg2hw.tag_1318.re;
  assign rcache_line[5][38].status_reg.status = reg2hw.status_1318.q;//status_reg_t'(reg2hw.status_1318.q);
  assign rcache_line[5][38].status_reg.qe    = reg2hw.status_1318.qe;
  assign rcache_line[5][38].status_reg.re    = reg2hw.status_1318.re;


  assign rcache_line[5][39].tag_reg.tag      = reg2hw.tag_1319.q;
  assign rcache_line[5][39].tag_reg.qe       = reg2hw.tag_1319.qe;
  assign rcache_line[5][39].tag_reg.re       = reg2hw.tag_1319.re;
  assign rcache_line[5][39].status_reg.status = reg2hw.status_1319.q;//status_reg_t'(reg2hw.status_1319.q);
  assign rcache_line[5][39].status_reg.qe    = reg2hw.status_1319.qe;
  assign rcache_line[5][39].status_reg.re    = reg2hw.status_1319.re;


  assign rcache_line[5][40].tag_reg.tag      = reg2hw.tag_1320.q;
  assign rcache_line[5][40].tag_reg.qe       = reg2hw.tag_1320.qe;
  assign rcache_line[5][40].tag_reg.re       = reg2hw.tag_1320.re;
  assign rcache_line[5][40].status_reg.status = reg2hw.status_1320.q;//status_reg_t'(reg2hw.status_1320.q);
  assign rcache_line[5][40].status_reg.qe    = reg2hw.status_1320.qe;
  assign rcache_line[5][40].status_reg.re    = reg2hw.status_1320.re;


  assign rcache_line[5][41].tag_reg.tag      = reg2hw.tag_1321.q;
  assign rcache_line[5][41].tag_reg.qe       = reg2hw.tag_1321.qe;
  assign rcache_line[5][41].tag_reg.re       = reg2hw.tag_1321.re;
  assign rcache_line[5][41].status_reg.status = reg2hw.status_1321.q;//status_reg_t'(reg2hw.status_1321.q);
  assign rcache_line[5][41].status_reg.qe    = reg2hw.status_1321.qe;
  assign rcache_line[5][41].status_reg.re    = reg2hw.status_1321.re;


  assign rcache_line[5][42].tag_reg.tag      = reg2hw.tag_1322.q;
  assign rcache_line[5][42].tag_reg.qe       = reg2hw.tag_1322.qe;
  assign rcache_line[5][42].tag_reg.re       = reg2hw.tag_1322.re;
  assign rcache_line[5][42].status_reg.status = reg2hw.status_1322.q;//status_reg_t'(reg2hw.status_1322.q);
  assign rcache_line[5][42].status_reg.qe    = reg2hw.status_1322.qe;
  assign rcache_line[5][42].status_reg.re    = reg2hw.status_1322.re;


  assign rcache_line[5][43].tag_reg.tag      = reg2hw.tag_1323.q;
  assign rcache_line[5][43].tag_reg.qe       = reg2hw.tag_1323.qe;
  assign rcache_line[5][43].tag_reg.re       = reg2hw.tag_1323.re;
  assign rcache_line[5][43].status_reg.status = reg2hw.status_1323.q;//status_reg_t'(reg2hw.status_1323.q);
  assign rcache_line[5][43].status_reg.qe    = reg2hw.status_1323.qe;
  assign rcache_line[5][43].status_reg.re    = reg2hw.status_1323.re;


  assign rcache_line[5][44].tag_reg.tag      = reg2hw.tag_1324.q;
  assign rcache_line[5][44].tag_reg.qe       = reg2hw.tag_1324.qe;
  assign rcache_line[5][44].tag_reg.re       = reg2hw.tag_1324.re;
  assign rcache_line[5][44].status_reg.status = reg2hw.status_1324.q;//status_reg_t'(reg2hw.status_1324.q);
  assign rcache_line[5][44].status_reg.qe    = reg2hw.status_1324.qe;
  assign rcache_line[5][44].status_reg.re    = reg2hw.status_1324.re;


  assign rcache_line[5][45].tag_reg.tag      = reg2hw.tag_1325.q;
  assign rcache_line[5][45].tag_reg.qe       = reg2hw.tag_1325.qe;
  assign rcache_line[5][45].tag_reg.re       = reg2hw.tag_1325.re;
  assign rcache_line[5][45].status_reg.status = reg2hw.status_1325.q;//status_reg_t'(reg2hw.status_1325.q);
  assign rcache_line[5][45].status_reg.qe    = reg2hw.status_1325.qe;
  assign rcache_line[5][45].status_reg.re    = reg2hw.status_1325.re;


  assign rcache_line[5][46].tag_reg.tag      = reg2hw.tag_1326.q;
  assign rcache_line[5][46].tag_reg.qe       = reg2hw.tag_1326.qe;
  assign rcache_line[5][46].tag_reg.re       = reg2hw.tag_1326.re;
  assign rcache_line[5][46].status_reg.status = reg2hw.status_1326.q;//status_reg_t'(reg2hw.status_1326.q);
  assign rcache_line[5][46].status_reg.qe    = reg2hw.status_1326.qe;
  assign rcache_line[5][46].status_reg.re    = reg2hw.status_1326.re;


  assign rcache_line[5][47].tag_reg.tag      = reg2hw.tag_1327.q;
  assign rcache_line[5][47].tag_reg.qe       = reg2hw.tag_1327.qe;
  assign rcache_line[5][47].tag_reg.re       = reg2hw.tag_1327.re;
  assign rcache_line[5][47].status_reg.status = reg2hw.status_1327.q;//status_reg_t'(reg2hw.status_1327.q);
  assign rcache_line[5][47].status_reg.qe    = reg2hw.status_1327.qe;
  assign rcache_line[5][47].status_reg.re    = reg2hw.status_1327.re;


  assign rcache_line[5][48].tag_reg.tag      = reg2hw.tag_1328.q;
  assign rcache_line[5][48].tag_reg.qe       = reg2hw.tag_1328.qe;
  assign rcache_line[5][48].tag_reg.re       = reg2hw.tag_1328.re;
  assign rcache_line[5][48].status_reg.status = reg2hw.status_1328.q;//status_reg_t'(reg2hw.status_1328.q);
  assign rcache_line[5][48].status_reg.qe    = reg2hw.status_1328.qe;
  assign rcache_line[5][48].status_reg.re    = reg2hw.status_1328.re;


  assign rcache_line[5][49].tag_reg.tag      = reg2hw.tag_1329.q;
  assign rcache_line[5][49].tag_reg.qe       = reg2hw.tag_1329.qe;
  assign rcache_line[5][49].tag_reg.re       = reg2hw.tag_1329.re;
  assign rcache_line[5][49].status_reg.status = reg2hw.status_1329.q;//status_reg_t'(reg2hw.status_1329.q);
  assign rcache_line[5][49].status_reg.qe    = reg2hw.status_1329.qe;
  assign rcache_line[5][49].status_reg.re    = reg2hw.status_1329.re;


  assign rcache_line[5][50].tag_reg.tag      = reg2hw.tag_1330.q;
  assign rcache_line[5][50].tag_reg.qe       = reg2hw.tag_1330.qe;
  assign rcache_line[5][50].tag_reg.re       = reg2hw.tag_1330.re;
  assign rcache_line[5][50].status_reg.status = reg2hw.status_1330.q;//status_reg_t'(reg2hw.status_1330.q);
  assign rcache_line[5][50].status_reg.qe    = reg2hw.status_1330.qe;
  assign rcache_line[5][50].status_reg.re    = reg2hw.status_1330.re;


  assign rcache_line[5][51].tag_reg.tag      = reg2hw.tag_1331.q;
  assign rcache_line[5][51].tag_reg.qe       = reg2hw.tag_1331.qe;
  assign rcache_line[5][51].tag_reg.re       = reg2hw.tag_1331.re;
  assign rcache_line[5][51].status_reg.status = reg2hw.status_1331.q;//status_reg_t'(reg2hw.status_1331.q);
  assign rcache_line[5][51].status_reg.qe    = reg2hw.status_1331.qe;
  assign rcache_line[5][51].status_reg.re    = reg2hw.status_1331.re;


  assign rcache_line[5][52].tag_reg.tag      = reg2hw.tag_1332.q;
  assign rcache_line[5][52].tag_reg.qe       = reg2hw.tag_1332.qe;
  assign rcache_line[5][52].tag_reg.re       = reg2hw.tag_1332.re;
  assign rcache_line[5][52].status_reg.status = reg2hw.status_1332.q;//status_reg_t'(reg2hw.status_1332.q);
  assign rcache_line[5][52].status_reg.qe    = reg2hw.status_1332.qe;
  assign rcache_line[5][52].status_reg.re    = reg2hw.status_1332.re;


  assign rcache_line[5][53].tag_reg.tag      = reg2hw.tag_1333.q;
  assign rcache_line[5][53].tag_reg.qe       = reg2hw.tag_1333.qe;
  assign rcache_line[5][53].tag_reg.re       = reg2hw.tag_1333.re;
  assign rcache_line[5][53].status_reg.status = reg2hw.status_1333.q;//status_reg_t'(reg2hw.status_1333.q);
  assign rcache_line[5][53].status_reg.qe    = reg2hw.status_1333.qe;
  assign rcache_line[5][53].status_reg.re    = reg2hw.status_1333.re;


  assign rcache_line[5][54].tag_reg.tag      = reg2hw.tag_1334.q;
  assign rcache_line[5][54].tag_reg.qe       = reg2hw.tag_1334.qe;
  assign rcache_line[5][54].tag_reg.re       = reg2hw.tag_1334.re;
  assign rcache_line[5][54].status_reg.status = reg2hw.status_1334.q;//status_reg_t'(reg2hw.status_1334.q);
  assign rcache_line[5][54].status_reg.qe    = reg2hw.status_1334.qe;
  assign rcache_line[5][54].status_reg.re    = reg2hw.status_1334.re;


  assign rcache_line[5][55].tag_reg.tag      = reg2hw.tag_1335.q;
  assign rcache_line[5][55].tag_reg.qe       = reg2hw.tag_1335.qe;
  assign rcache_line[5][55].tag_reg.re       = reg2hw.tag_1335.re;
  assign rcache_line[5][55].status_reg.status = reg2hw.status_1335.q;//status_reg_t'(reg2hw.status_1335.q);
  assign rcache_line[5][55].status_reg.qe    = reg2hw.status_1335.qe;
  assign rcache_line[5][55].status_reg.re    = reg2hw.status_1335.re;


  assign rcache_line[5][56].tag_reg.tag      = reg2hw.tag_1336.q;
  assign rcache_line[5][56].tag_reg.qe       = reg2hw.tag_1336.qe;
  assign rcache_line[5][56].tag_reg.re       = reg2hw.tag_1336.re;
  assign rcache_line[5][56].status_reg.status = reg2hw.status_1336.q;//status_reg_t'(reg2hw.status_1336.q);
  assign rcache_line[5][56].status_reg.qe    = reg2hw.status_1336.qe;
  assign rcache_line[5][56].status_reg.re    = reg2hw.status_1336.re;


  assign rcache_line[5][57].tag_reg.tag      = reg2hw.tag_1337.q;
  assign rcache_line[5][57].tag_reg.qe       = reg2hw.tag_1337.qe;
  assign rcache_line[5][57].tag_reg.re       = reg2hw.tag_1337.re;
  assign rcache_line[5][57].status_reg.status = reg2hw.status_1337.q;//status_reg_t'(reg2hw.status_1337.q);
  assign rcache_line[5][57].status_reg.qe    = reg2hw.status_1337.qe;
  assign rcache_line[5][57].status_reg.re    = reg2hw.status_1337.re;


  assign rcache_line[5][58].tag_reg.tag      = reg2hw.tag_1338.q;
  assign rcache_line[5][58].tag_reg.qe       = reg2hw.tag_1338.qe;
  assign rcache_line[5][58].tag_reg.re       = reg2hw.tag_1338.re;
  assign rcache_line[5][58].status_reg.status = reg2hw.status_1338.q;//status_reg_t'(reg2hw.status_1338.q);
  assign rcache_line[5][58].status_reg.qe    = reg2hw.status_1338.qe;
  assign rcache_line[5][58].status_reg.re    = reg2hw.status_1338.re;


  assign rcache_line[5][59].tag_reg.tag      = reg2hw.tag_1339.q;
  assign rcache_line[5][59].tag_reg.qe       = reg2hw.tag_1339.qe;
  assign rcache_line[5][59].tag_reg.re       = reg2hw.tag_1339.re;
  assign rcache_line[5][59].status_reg.status = reg2hw.status_1339.q;//status_reg_t'(reg2hw.status_1339.q);
  assign rcache_line[5][59].status_reg.qe    = reg2hw.status_1339.qe;
  assign rcache_line[5][59].status_reg.re    = reg2hw.status_1339.re;


  assign rcache_line[5][60].tag_reg.tag      = reg2hw.tag_1340.q;
  assign rcache_line[5][60].tag_reg.qe       = reg2hw.tag_1340.qe;
  assign rcache_line[5][60].tag_reg.re       = reg2hw.tag_1340.re;
  assign rcache_line[5][60].status_reg.status = reg2hw.status_1340.q;//status_reg_t'(reg2hw.status_1340.q);
  assign rcache_line[5][60].status_reg.qe    = reg2hw.status_1340.qe;
  assign rcache_line[5][60].status_reg.re    = reg2hw.status_1340.re;


  assign rcache_line[5][61].tag_reg.tag      = reg2hw.tag_1341.q;
  assign rcache_line[5][61].tag_reg.qe       = reg2hw.tag_1341.qe;
  assign rcache_line[5][61].tag_reg.re       = reg2hw.tag_1341.re;
  assign rcache_line[5][61].status_reg.status = reg2hw.status_1341.q;//status_reg_t'(reg2hw.status_1341.q);
  assign rcache_line[5][61].status_reg.qe    = reg2hw.status_1341.qe;
  assign rcache_line[5][61].status_reg.re    = reg2hw.status_1341.re;


  assign rcache_line[5][62].tag_reg.tag      = reg2hw.tag_1342.q;
  assign rcache_line[5][62].tag_reg.qe       = reg2hw.tag_1342.qe;
  assign rcache_line[5][62].tag_reg.re       = reg2hw.tag_1342.re;
  assign rcache_line[5][62].status_reg.status = reg2hw.status_1342.q;//status_reg_t'(reg2hw.status_1342.q);
  assign rcache_line[5][62].status_reg.qe    = reg2hw.status_1342.qe;
  assign rcache_line[5][62].status_reg.re    = reg2hw.status_1342.re;


  assign rcache_line[5][63].tag_reg.tag      = reg2hw.tag_1343.q;
  assign rcache_line[5][63].tag_reg.qe       = reg2hw.tag_1343.qe;
  assign rcache_line[5][63].tag_reg.re       = reg2hw.tag_1343.re;
  assign rcache_line[5][63].status_reg.status = reg2hw.status_1343.q;//status_reg_t'(reg2hw.status_1343.q);
  assign rcache_line[5][63].status_reg.qe    = reg2hw.status_1343.qe;
  assign rcache_line[5][63].status_reg.re    = reg2hw.status_1343.re;


  assign rcache_line[5][64].tag_reg.tag      = reg2hw.tag_1344.q;
  assign rcache_line[5][64].tag_reg.qe       = reg2hw.tag_1344.qe;
  assign rcache_line[5][64].tag_reg.re       = reg2hw.tag_1344.re;
  assign rcache_line[5][64].status_reg.status = reg2hw.status_1344.q;//status_reg_t'(reg2hw.status_1344.q);
  assign rcache_line[5][64].status_reg.qe    = reg2hw.status_1344.qe;
  assign rcache_line[5][64].status_reg.re    = reg2hw.status_1344.re;


  assign rcache_line[5][65].tag_reg.tag      = reg2hw.tag_1345.q;
  assign rcache_line[5][65].tag_reg.qe       = reg2hw.tag_1345.qe;
  assign rcache_line[5][65].tag_reg.re       = reg2hw.tag_1345.re;
  assign rcache_line[5][65].status_reg.status = reg2hw.status_1345.q;//status_reg_t'(reg2hw.status_1345.q);
  assign rcache_line[5][65].status_reg.qe    = reg2hw.status_1345.qe;
  assign rcache_line[5][65].status_reg.re    = reg2hw.status_1345.re;


  assign rcache_line[5][66].tag_reg.tag      = reg2hw.tag_1346.q;
  assign rcache_line[5][66].tag_reg.qe       = reg2hw.tag_1346.qe;
  assign rcache_line[5][66].tag_reg.re       = reg2hw.tag_1346.re;
  assign rcache_line[5][66].status_reg.status = reg2hw.status_1346.q;//status_reg_t'(reg2hw.status_1346.q);
  assign rcache_line[5][66].status_reg.qe    = reg2hw.status_1346.qe;
  assign rcache_line[5][66].status_reg.re    = reg2hw.status_1346.re;


  assign rcache_line[5][67].tag_reg.tag      = reg2hw.tag_1347.q;
  assign rcache_line[5][67].tag_reg.qe       = reg2hw.tag_1347.qe;
  assign rcache_line[5][67].tag_reg.re       = reg2hw.tag_1347.re;
  assign rcache_line[5][67].status_reg.status = reg2hw.status_1347.q;//status_reg_t'(reg2hw.status_1347.q);
  assign rcache_line[5][67].status_reg.qe    = reg2hw.status_1347.qe;
  assign rcache_line[5][67].status_reg.re    = reg2hw.status_1347.re;


  assign rcache_line[5][68].tag_reg.tag      = reg2hw.tag_1348.q;
  assign rcache_line[5][68].tag_reg.qe       = reg2hw.tag_1348.qe;
  assign rcache_line[5][68].tag_reg.re       = reg2hw.tag_1348.re;
  assign rcache_line[5][68].status_reg.status = reg2hw.status_1348.q;//status_reg_t'(reg2hw.status_1348.q);
  assign rcache_line[5][68].status_reg.qe    = reg2hw.status_1348.qe;
  assign rcache_line[5][68].status_reg.re    = reg2hw.status_1348.re;


  assign rcache_line[5][69].tag_reg.tag      = reg2hw.tag_1349.q;
  assign rcache_line[5][69].tag_reg.qe       = reg2hw.tag_1349.qe;
  assign rcache_line[5][69].tag_reg.re       = reg2hw.tag_1349.re;
  assign rcache_line[5][69].status_reg.status = reg2hw.status_1349.q;//status_reg_t'(reg2hw.status_1349.q);
  assign rcache_line[5][69].status_reg.qe    = reg2hw.status_1349.qe;
  assign rcache_line[5][69].status_reg.re    = reg2hw.status_1349.re;


  assign rcache_line[5][70].tag_reg.tag      = reg2hw.tag_1350.q;
  assign rcache_line[5][70].tag_reg.qe       = reg2hw.tag_1350.qe;
  assign rcache_line[5][70].tag_reg.re       = reg2hw.tag_1350.re;
  assign rcache_line[5][70].status_reg.status = reg2hw.status_1350.q;//status_reg_t'(reg2hw.status_1350.q);
  assign rcache_line[5][70].status_reg.qe    = reg2hw.status_1350.qe;
  assign rcache_line[5][70].status_reg.re    = reg2hw.status_1350.re;


  assign rcache_line[5][71].tag_reg.tag      = reg2hw.tag_1351.q;
  assign rcache_line[5][71].tag_reg.qe       = reg2hw.tag_1351.qe;
  assign rcache_line[5][71].tag_reg.re       = reg2hw.tag_1351.re;
  assign rcache_line[5][71].status_reg.status = reg2hw.status_1351.q;//status_reg_t'(reg2hw.status_1351.q);
  assign rcache_line[5][71].status_reg.qe    = reg2hw.status_1351.qe;
  assign rcache_line[5][71].status_reg.re    = reg2hw.status_1351.re;


  assign rcache_line[5][72].tag_reg.tag      = reg2hw.tag_1352.q;
  assign rcache_line[5][72].tag_reg.qe       = reg2hw.tag_1352.qe;
  assign rcache_line[5][72].tag_reg.re       = reg2hw.tag_1352.re;
  assign rcache_line[5][72].status_reg.status = reg2hw.status_1352.q;//status_reg_t'(reg2hw.status_1352.q);
  assign rcache_line[5][72].status_reg.qe    = reg2hw.status_1352.qe;
  assign rcache_line[5][72].status_reg.re    = reg2hw.status_1352.re;


  assign rcache_line[5][73].tag_reg.tag      = reg2hw.tag_1353.q;
  assign rcache_line[5][73].tag_reg.qe       = reg2hw.tag_1353.qe;
  assign rcache_line[5][73].tag_reg.re       = reg2hw.tag_1353.re;
  assign rcache_line[5][73].status_reg.status = reg2hw.status_1353.q;//status_reg_t'(reg2hw.status_1353.q);
  assign rcache_line[5][73].status_reg.qe    = reg2hw.status_1353.qe;
  assign rcache_line[5][73].status_reg.re    = reg2hw.status_1353.re;


  assign rcache_line[5][74].tag_reg.tag      = reg2hw.tag_1354.q;
  assign rcache_line[5][74].tag_reg.qe       = reg2hw.tag_1354.qe;
  assign rcache_line[5][74].tag_reg.re       = reg2hw.tag_1354.re;
  assign rcache_line[5][74].status_reg.status = reg2hw.status_1354.q;//status_reg_t'(reg2hw.status_1354.q);
  assign rcache_line[5][74].status_reg.qe    = reg2hw.status_1354.qe;
  assign rcache_line[5][74].status_reg.re    = reg2hw.status_1354.re;


  assign rcache_line[5][75].tag_reg.tag      = reg2hw.tag_1355.q;
  assign rcache_line[5][75].tag_reg.qe       = reg2hw.tag_1355.qe;
  assign rcache_line[5][75].tag_reg.re       = reg2hw.tag_1355.re;
  assign rcache_line[5][75].status_reg.status = reg2hw.status_1355.q;//status_reg_t'(reg2hw.status_1355.q);
  assign rcache_line[5][75].status_reg.qe    = reg2hw.status_1355.qe;
  assign rcache_line[5][75].status_reg.re    = reg2hw.status_1355.re;


  assign rcache_line[5][76].tag_reg.tag      = reg2hw.tag_1356.q;
  assign rcache_line[5][76].tag_reg.qe       = reg2hw.tag_1356.qe;
  assign rcache_line[5][76].tag_reg.re       = reg2hw.tag_1356.re;
  assign rcache_line[5][76].status_reg.status = reg2hw.status_1356.q;//status_reg_t'(reg2hw.status_1356.q);
  assign rcache_line[5][76].status_reg.qe    = reg2hw.status_1356.qe;
  assign rcache_line[5][76].status_reg.re    = reg2hw.status_1356.re;


  assign rcache_line[5][77].tag_reg.tag      = reg2hw.tag_1357.q;
  assign rcache_line[5][77].tag_reg.qe       = reg2hw.tag_1357.qe;
  assign rcache_line[5][77].tag_reg.re       = reg2hw.tag_1357.re;
  assign rcache_line[5][77].status_reg.status = reg2hw.status_1357.q;//status_reg_t'(reg2hw.status_1357.q);
  assign rcache_line[5][77].status_reg.qe    = reg2hw.status_1357.qe;
  assign rcache_line[5][77].status_reg.re    = reg2hw.status_1357.re;


  assign rcache_line[5][78].tag_reg.tag      = reg2hw.tag_1358.q;
  assign rcache_line[5][78].tag_reg.qe       = reg2hw.tag_1358.qe;
  assign rcache_line[5][78].tag_reg.re       = reg2hw.tag_1358.re;
  assign rcache_line[5][78].status_reg.status = reg2hw.status_1358.q;//status_reg_t'(reg2hw.status_1358.q);
  assign rcache_line[5][78].status_reg.qe    = reg2hw.status_1358.qe;
  assign rcache_line[5][78].status_reg.re    = reg2hw.status_1358.re;


  assign rcache_line[5][79].tag_reg.tag      = reg2hw.tag_1359.q;
  assign rcache_line[5][79].tag_reg.qe       = reg2hw.tag_1359.qe;
  assign rcache_line[5][79].tag_reg.re       = reg2hw.tag_1359.re;
  assign rcache_line[5][79].status_reg.status = reg2hw.status_1359.q;//status_reg_t'(reg2hw.status_1359.q);
  assign rcache_line[5][79].status_reg.qe    = reg2hw.status_1359.qe;
  assign rcache_line[5][79].status_reg.re    = reg2hw.status_1359.re;


  assign rcache_line[5][80].tag_reg.tag      = reg2hw.tag_1360.q;
  assign rcache_line[5][80].tag_reg.qe       = reg2hw.tag_1360.qe;
  assign rcache_line[5][80].tag_reg.re       = reg2hw.tag_1360.re;
  assign rcache_line[5][80].status_reg.status = reg2hw.status_1360.q;//status_reg_t'(reg2hw.status_1360.q);
  assign rcache_line[5][80].status_reg.qe    = reg2hw.status_1360.qe;
  assign rcache_line[5][80].status_reg.re    = reg2hw.status_1360.re;


  assign rcache_line[5][81].tag_reg.tag      = reg2hw.tag_1361.q;
  assign rcache_line[5][81].tag_reg.qe       = reg2hw.tag_1361.qe;
  assign rcache_line[5][81].tag_reg.re       = reg2hw.tag_1361.re;
  assign rcache_line[5][81].status_reg.status = reg2hw.status_1361.q;//status_reg_t'(reg2hw.status_1361.q);
  assign rcache_line[5][81].status_reg.qe    = reg2hw.status_1361.qe;
  assign rcache_line[5][81].status_reg.re    = reg2hw.status_1361.re;


  assign rcache_line[5][82].tag_reg.tag      = reg2hw.tag_1362.q;
  assign rcache_line[5][82].tag_reg.qe       = reg2hw.tag_1362.qe;
  assign rcache_line[5][82].tag_reg.re       = reg2hw.tag_1362.re;
  assign rcache_line[5][82].status_reg.status = reg2hw.status_1362.q;//status_reg_t'(reg2hw.status_1362.q);
  assign rcache_line[5][82].status_reg.qe    = reg2hw.status_1362.qe;
  assign rcache_line[5][82].status_reg.re    = reg2hw.status_1362.re;


  assign rcache_line[5][83].tag_reg.tag      = reg2hw.tag_1363.q;
  assign rcache_line[5][83].tag_reg.qe       = reg2hw.tag_1363.qe;
  assign rcache_line[5][83].tag_reg.re       = reg2hw.tag_1363.re;
  assign rcache_line[5][83].status_reg.status = reg2hw.status_1363.q;//status_reg_t'(reg2hw.status_1363.q);
  assign rcache_line[5][83].status_reg.qe    = reg2hw.status_1363.qe;
  assign rcache_line[5][83].status_reg.re    = reg2hw.status_1363.re;


  assign rcache_line[5][84].tag_reg.tag      = reg2hw.tag_1364.q;
  assign rcache_line[5][84].tag_reg.qe       = reg2hw.tag_1364.qe;
  assign rcache_line[5][84].tag_reg.re       = reg2hw.tag_1364.re;
  assign rcache_line[5][84].status_reg.status = reg2hw.status_1364.q;//status_reg_t'(reg2hw.status_1364.q);
  assign rcache_line[5][84].status_reg.qe    = reg2hw.status_1364.qe;
  assign rcache_line[5][84].status_reg.re    = reg2hw.status_1364.re;


  assign rcache_line[5][85].tag_reg.tag      = reg2hw.tag_1365.q;
  assign rcache_line[5][85].tag_reg.qe       = reg2hw.tag_1365.qe;
  assign rcache_line[5][85].tag_reg.re       = reg2hw.tag_1365.re;
  assign rcache_line[5][85].status_reg.status = reg2hw.status_1365.q;//status_reg_t'(reg2hw.status_1365.q);
  assign rcache_line[5][85].status_reg.qe    = reg2hw.status_1365.qe;
  assign rcache_line[5][85].status_reg.re    = reg2hw.status_1365.re;


  assign rcache_line[5][86].tag_reg.tag      = reg2hw.tag_1366.q;
  assign rcache_line[5][86].tag_reg.qe       = reg2hw.tag_1366.qe;
  assign rcache_line[5][86].tag_reg.re       = reg2hw.tag_1366.re;
  assign rcache_line[5][86].status_reg.status = reg2hw.status_1366.q;//status_reg_t'(reg2hw.status_1366.q);
  assign rcache_line[5][86].status_reg.qe    = reg2hw.status_1366.qe;
  assign rcache_line[5][86].status_reg.re    = reg2hw.status_1366.re;


  assign rcache_line[5][87].tag_reg.tag      = reg2hw.tag_1367.q;
  assign rcache_line[5][87].tag_reg.qe       = reg2hw.tag_1367.qe;
  assign rcache_line[5][87].tag_reg.re       = reg2hw.tag_1367.re;
  assign rcache_line[5][87].status_reg.status = reg2hw.status_1367.q;//status_reg_t'(reg2hw.status_1367.q);
  assign rcache_line[5][87].status_reg.qe    = reg2hw.status_1367.qe;
  assign rcache_line[5][87].status_reg.re    = reg2hw.status_1367.re;


  assign rcache_line[5][88].tag_reg.tag      = reg2hw.tag_1368.q;
  assign rcache_line[5][88].tag_reg.qe       = reg2hw.tag_1368.qe;
  assign rcache_line[5][88].tag_reg.re       = reg2hw.tag_1368.re;
  assign rcache_line[5][88].status_reg.status = reg2hw.status_1368.q;//status_reg_t'(reg2hw.status_1368.q);
  assign rcache_line[5][88].status_reg.qe    = reg2hw.status_1368.qe;
  assign rcache_line[5][88].status_reg.re    = reg2hw.status_1368.re;


  assign rcache_line[5][89].tag_reg.tag      = reg2hw.tag_1369.q;
  assign rcache_line[5][89].tag_reg.qe       = reg2hw.tag_1369.qe;
  assign rcache_line[5][89].tag_reg.re       = reg2hw.tag_1369.re;
  assign rcache_line[5][89].status_reg.status = reg2hw.status_1369.q;//status_reg_t'(reg2hw.status_1369.q);
  assign rcache_line[5][89].status_reg.qe    = reg2hw.status_1369.qe;
  assign rcache_line[5][89].status_reg.re    = reg2hw.status_1369.re;


  assign rcache_line[5][90].tag_reg.tag      = reg2hw.tag_1370.q;
  assign rcache_line[5][90].tag_reg.qe       = reg2hw.tag_1370.qe;
  assign rcache_line[5][90].tag_reg.re       = reg2hw.tag_1370.re;
  assign rcache_line[5][90].status_reg.status = reg2hw.status_1370.q;//status_reg_t'(reg2hw.status_1370.q);
  assign rcache_line[5][90].status_reg.qe    = reg2hw.status_1370.qe;
  assign rcache_line[5][90].status_reg.re    = reg2hw.status_1370.re;


  assign rcache_line[5][91].tag_reg.tag      = reg2hw.tag_1371.q;
  assign rcache_line[5][91].tag_reg.qe       = reg2hw.tag_1371.qe;
  assign rcache_line[5][91].tag_reg.re       = reg2hw.tag_1371.re;
  assign rcache_line[5][91].status_reg.status = reg2hw.status_1371.q;//status_reg_t'(reg2hw.status_1371.q);
  assign rcache_line[5][91].status_reg.qe    = reg2hw.status_1371.qe;
  assign rcache_line[5][91].status_reg.re    = reg2hw.status_1371.re;


  assign rcache_line[5][92].tag_reg.tag      = reg2hw.tag_1372.q;
  assign rcache_line[5][92].tag_reg.qe       = reg2hw.tag_1372.qe;
  assign rcache_line[5][92].tag_reg.re       = reg2hw.tag_1372.re;
  assign rcache_line[5][92].status_reg.status = reg2hw.status_1372.q;//status_reg_t'(reg2hw.status_1372.q);
  assign rcache_line[5][92].status_reg.qe    = reg2hw.status_1372.qe;
  assign rcache_line[5][92].status_reg.re    = reg2hw.status_1372.re;


  assign rcache_line[5][93].tag_reg.tag      = reg2hw.tag_1373.q;
  assign rcache_line[5][93].tag_reg.qe       = reg2hw.tag_1373.qe;
  assign rcache_line[5][93].tag_reg.re       = reg2hw.tag_1373.re;
  assign rcache_line[5][93].status_reg.status = reg2hw.status_1373.q;//status_reg_t'(reg2hw.status_1373.q);
  assign rcache_line[5][93].status_reg.qe    = reg2hw.status_1373.qe;
  assign rcache_line[5][93].status_reg.re    = reg2hw.status_1373.re;


  assign rcache_line[5][94].tag_reg.tag      = reg2hw.tag_1374.q;
  assign rcache_line[5][94].tag_reg.qe       = reg2hw.tag_1374.qe;
  assign rcache_line[5][94].tag_reg.re       = reg2hw.tag_1374.re;
  assign rcache_line[5][94].status_reg.status = reg2hw.status_1374.q;//status_reg_t'(reg2hw.status_1374.q);
  assign rcache_line[5][94].status_reg.qe    = reg2hw.status_1374.qe;
  assign rcache_line[5][94].status_reg.re    = reg2hw.status_1374.re;


  assign rcache_line[5][95].tag_reg.tag      = reg2hw.tag_1375.q;
  assign rcache_line[5][95].tag_reg.qe       = reg2hw.tag_1375.qe;
  assign rcache_line[5][95].tag_reg.re       = reg2hw.tag_1375.re;
  assign rcache_line[5][95].status_reg.status = reg2hw.status_1375.q;//status_reg_t'(reg2hw.status_1375.q);
  assign rcache_line[5][95].status_reg.qe    = reg2hw.status_1375.qe;
  assign rcache_line[5][95].status_reg.re    = reg2hw.status_1375.re;


  assign rcache_line[5][96].tag_reg.tag      = reg2hw.tag_1376.q;
  assign rcache_line[5][96].tag_reg.qe       = reg2hw.tag_1376.qe;
  assign rcache_line[5][96].tag_reg.re       = reg2hw.tag_1376.re;
  assign rcache_line[5][96].status_reg.status = reg2hw.status_1376.q;//status_reg_t'(reg2hw.status_1376.q);
  assign rcache_line[5][96].status_reg.qe    = reg2hw.status_1376.qe;
  assign rcache_line[5][96].status_reg.re    = reg2hw.status_1376.re;


  assign rcache_line[5][97].tag_reg.tag      = reg2hw.tag_1377.q;
  assign rcache_line[5][97].tag_reg.qe       = reg2hw.tag_1377.qe;
  assign rcache_line[5][97].tag_reg.re       = reg2hw.tag_1377.re;
  assign rcache_line[5][97].status_reg.status = reg2hw.status_1377.q;//status_reg_t'(reg2hw.status_1377.q);
  assign rcache_line[5][97].status_reg.qe    = reg2hw.status_1377.qe;
  assign rcache_line[5][97].status_reg.re    = reg2hw.status_1377.re;


  assign rcache_line[5][98].tag_reg.tag      = reg2hw.tag_1378.q;
  assign rcache_line[5][98].tag_reg.qe       = reg2hw.tag_1378.qe;
  assign rcache_line[5][98].tag_reg.re       = reg2hw.tag_1378.re;
  assign rcache_line[5][98].status_reg.status = reg2hw.status_1378.q;//status_reg_t'(reg2hw.status_1378.q);
  assign rcache_line[5][98].status_reg.qe    = reg2hw.status_1378.qe;
  assign rcache_line[5][98].status_reg.re    = reg2hw.status_1378.re;


  assign rcache_line[5][99].tag_reg.tag      = reg2hw.tag_1379.q;
  assign rcache_line[5][99].tag_reg.qe       = reg2hw.tag_1379.qe;
  assign rcache_line[5][99].tag_reg.re       = reg2hw.tag_1379.re;
  assign rcache_line[5][99].status_reg.status = reg2hw.status_1379.q;//status_reg_t'(reg2hw.status_1379.q);
  assign rcache_line[5][99].status_reg.qe    = reg2hw.status_1379.qe;
  assign rcache_line[5][99].status_reg.re    = reg2hw.status_1379.re;


  assign rcache_line[5][100].tag_reg.tag      = reg2hw.tag_1380.q;
  assign rcache_line[5][100].tag_reg.qe       = reg2hw.tag_1380.qe;
  assign rcache_line[5][100].tag_reg.re       = reg2hw.tag_1380.re;
  assign rcache_line[5][100].status_reg.status = reg2hw.status_1380.q;//status_reg_t'(reg2hw.status_1380.q);
  assign rcache_line[5][100].status_reg.qe    = reg2hw.status_1380.qe;
  assign rcache_line[5][100].status_reg.re    = reg2hw.status_1380.re;


  assign rcache_line[5][101].tag_reg.tag      = reg2hw.tag_1381.q;
  assign rcache_line[5][101].tag_reg.qe       = reg2hw.tag_1381.qe;
  assign rcache_line[5][101].tag_reg.re       = reg2hw.tag_1381.re;
  assign rcache_line[5][101].status_reg.status = reg2hw.status_1381.q;//status_reg_t'(reg2hw.status_1381.q);
  assign rcache_line[5][101].status_reg.qe    = reg2hw.status_1381.qe;
  assign rcache_line[5][101].status_reg.re    = reg2hw.status_1381.re;


  assign rcache_line[5][102].tag_reg.tag      = reg2hw.tag_1382.q;
  assign rcache_line[5][102].tag_reg.qe       = reg2hw.tag_1382.qe;
  assign rcache_line[5][102].tag_reg.re       = reg2hw.tag_1382.re;
  assign rcache_line[5][102].status_reg.status = reg2hw.status_1382.q;//status_reg_t'(reg2hw.status_1382.q);
  assign rcache_line[5][102].status_reg.qe    = reg2hw.status_1382.qe;
  assign rcache_line[5][102].status_reg.re    = reg2hw.status_1382.re;


  assign rcache_line[5][103].tag_reg.tag      = reg2hw.tag_1383.q;
  assign rcache_line[5][103].tag_reg.qe       = reg2hw.tag_1383.qe;
  assign rcache_line[5][103].tag_reg.re       = reg2hw.tag_1383.re;
  assign rcache_line[5][103].status_reg.status = reg2hw.status_1383.q;//status_reg_t'(reg2hw.status_1383.q);
  assign rcache_line[5][103].status_reg.qe    = reg2hw.status_1383.qe;
  assign rcache_line[5][103].status_reg.re    = reg2hw.status_1383.re;


  assign rcache_line[5][104].tag_reg.tag      = reg2hw.tag_1384.q;
  assign rcache_line[5][104].tag_reg.qe       = reg2hw.tag_1384.qe;
  assign rcache_line[5][104].tag_reg.re       = reg2hw.tag_1384.re;
  assign rcache_line[5][104].status_reg.status = reg2hw.status_1384.q;//status_reg_t'(reg2hw.status_1384.q);
  assign rcache_line[5][104].status_reg.qe    = reg2hw.status_1384.qe;
  assign rcache_line[5][104].status_reg.re    = reg2hw.status_1384.re;


  assign rcache_line[5][105].tag_reg.tag      = reg2hw.tag_1385.q;
  assign rcache_line[5][105].tag_reg.qe       = reg2hw.tag_1385.qe;
  assign rcache_line[5][105].tag_reg.re       = reg2hw.tag_1385.re;
  assign rcache_line[5][105].status_reg.status = reg2hw.status_1385.q;//status_reg_t'(reg2hw.status_1385.q);
  assign rcache_line[5][105].status_reg.qe    = reg2hw.status_1385.qe;
  assign rcache_line[5][105].status_reg.re    = reg2hw.status_1385.re;


  assign rcache_line[5][106].tag_reg.tag      = reg2hw.tag_1386.q;
  assign rcache_line[5][106].tag_reg.qe       = reg2hw.tag_1386.qe;
  assign rcache_line[5][106].tag_reg.re       = reg2hw.tag_1386.re;
  assign rcache_line[5][106].status_reg.status = reg2hw.status_1386.q;//status_reg_t'(reg2hw.status_1386.q);
  assign rcache_line[5][106].status_reg.qe    = reg2hw.status_1386.qe;
  assign rcache_line[5][106].status_reg.re    = reg2hw.status_1386.re;


  assign rcache_line[5][107].tag_reg.tag      = reg2hw.tag_1387.q;
  assign rcache_line[5][107].tag_reg.qe       = reg2hw.tag_1387.qe;
  assign rcache_line[5][107].tag_reg.re       = reg2hw.tag_1387.re;
  assign rcache_line[5][107].status_reg.status = reg2hw.status_1387.q;//status_reg_t'(reg2hw.status_1387.q);
  assign rcache_line[5][107].status_reg.qe    = reg2hw.status_1387.qe;
  assign rcache_line[5][107].status_reg.re    = reg2hw.status_1387.re;


  assign rcache_line[5][108].tag_reg.tag      = reg2hw.tag_1388.q;
  assign rcache_line[5][108].tag_reg.qe       = reg2hw.tag_1388.qe;
  assign rcache_line[5][108].tag_reg.re       = reg2hw.tag_1388.re;
  assign rcache_line[5][108].status_reg.status = reg2hw.status_1388.q;//status_reg_t'(reg2hw.status_1388.q);
  assign rcache_line[5][108].status_reg.qe    = reg2hw.status_1388.qe;
  assign rcache_line[5][108].status_reg.re    = reg2hw.status_1388.re;


  assign rcache_line[5][109].tag_reg.tag      = reg2hw.tag_1389.q;
  assign rcache_line[5][109].tag_reg.qe       = reg2hw.tag_1389.qe;
  assign rcache_line[5][109].tag_reg.re       = reg2hw.tag_1389.re;
  assign rcache_line[5][109].status_reg.status = reg2hw.status_1389.q;//status_reg_t'(reg2hw.status_1389.q);
  assign rcache_line[5][109].status_reg.qe    = reg2hw.status_1389.qe;
  assign rcache_line[5][109].status_reg.re    = reg2hw.status_1389.re;


  assign rcache_line[5][110].tag_reg.tag      = reg2hw.tag_1390.q;
  assign rcache_line[5][110].tag_reg.qe       = reg2hw.tag_1390.qe;
  assign rcache_line[5][110].tag_reg.re       = reg2hw.tag_1390.re;
  assign rcache_line[5][110].status_reg.status = reg2hw.status_1390.q;//status_reg_t'(reg2hw.status_1390.q);
  assign rcache_line[5][110].status_reg.qe    = reg2hw.status_1390.qe;
  assign rcache_line[5][110].status_reg.re    = reg2hw.status_1390.re;


  assign rcache_line[5][111].tag_reg.tag      = reg2hw.tag_1391.q;
  assign rcache_line[5][111].tag_reg.qe       = reg2hw.tag_1391.qe;
  assign rcache_line[5][111].tag_reg.re       = reg2hw.tag_1391.re;
  assign rcache_line[5][111].status_reg.status = reg2hw.status_1391.q;//status_reg_t'(reg2hw.status_1391.q);
  assign rcache_line[5][111].status_reg.qe    = reg2hw.status_1391.qe;
  assign rcache_line[5][111].status_reg.re    = reg2hw.status_1391.re;


  assign rcache_line[5][112].tag_reg.tag      = reg2hw.tag_1392.q;
  assign rcache_line[5][112].tag_reg.qe       = reg2hw.tag_1392.qe;
  assign rcache_line[5][112].tag_reg.re       = reg2hw.tag_1392.re;
  assign rcache_line[5][112].status_reg.status = reg2hw.status_1392.q;//status_reg_t'(reg2hw.status_1392.q);
  assign rcache_line[5][112].status_reg.qe    = reg2hw.status_1392.qe;
  assign rcache_line[5][112].status_reg.re    = reg2hw.status_1392.re;


  assign rcache_line[5][113].tag_reg.tag      = reg2hw.tag_1393.q;
  assign rcache_line[5][113].tag_reg.qe       = reg2hw.tag_1393.qe;
  assign rcache_line[5][113].tag_reg.re       = reg2hw.tag_1393.re;
  assign rcache_line[5][113].status_reg.status = reg2hw.status_1393.q;//status_reg_t'(reg2hw.status_1393.q);
  assign rcache_line[5][113].status_reg.qe    = reg2hw.status_1393.qe;
  assign rcache_line[5][113].status_reg.re    = reg2hw.status_1393.re;


  assign rcache_line[5][114].tag_reg.tag      = reg2hw.tag_1394.q;
  assign rcache_line[5][114].tag_reg.qe       = reg2hw.tag_1394.qe;
  assign rcache_line[5][114].tag_reg.re       = reg2hw.tag_1394.re;
  assign rcache_line[5][114].status_reg.status = reg2hw.status_1394.q;//status_reg_t'(reg2hw.status_1394.q);
  assign rcache_line[5][114].status_reg.qe    = reg2hw.status_1394.qe;
  assign rcache_line[5][114].status_reg.re    = reg2hw.status_1394.re;


  assign rcache_line[5][115].tag_reg.tag      = reg2hw.tag_1395.q;
  assign rcache_line[5][115].tag_reg.qe       = reg2hw.tag_1395.qe;
  assign rcache_line[5][115].tag_reg.re       = reg2hw.tag_1395.re;
  assign rcache_line[5][115].status_reg.status = reg2hw.status_1395.q;//status_reg_t'(reg2hw.status_1395.q);
  assign rcache_line[5][115].status_reg.qe    = reg2hw.status_1395.qe;
  assign rcache_line[5][115].status_reg.re    = reg2hw.status_1395.re;


  assign rcache_line[5][116].tag_reg.tag      = reg2hw.tag_1396.q;
  assign rcache_line[5][116].tag_reg.qe       = reg2hw.tag_1396.qe;
  assign rcache_line[5][116].tag_reg.re       = reg2hw.tag_1396.re;
  assign rcache_line[5][116].status_reg.status = reg2hw.status_1396.q;//status_reg_t'(reg2hw.status_1396.q);
  assign rcache_line[5][116].status_reg.qe    = reg2hw.status_1396.qe;
  assign rcache_line[5][116].status_reg.re    = reg2hw.status_1396.re;


  assign rcache_line[5][117].tag_reg.tag      = reg2hw.tag_1397.q;
  assign rcache_line[5][117].tag_reg.qe       = reg2hw.tag_1397.qe;
  assign rcache_line[5][117].tag_reg.re       = reg2hw.tag_1397.re;
  assign rcache_line[5][117].status_reg.status = reg2hw.status_1397.q;//status_reg_t'(reg2hw.status_1397.q);
  assign rcache_line[5][117].status_reg.qe    = reg2hw.status_1397.qe;
  assign rcache_line[5][117].status_reg.re    = reg2hw.status_1397.re;


  assign rcache_line[5][118].tag_reg.tag      = reg2hw.tag_1398.q;
  assign rcache_line[5][118].tag_reg.qe       = reg2hw.tag_1398.qe;
  assign rcache_line[5][118].tag_reg.re       = reg2hw.tag_1398.re;
  assign rcache_line[5][118].status_reg.status = reg2hw.status_1398.q;//status_reg_t'(reg2hw.status_1398.q);
  assign rcache_line[5][118].status_reg.qe    = reg2hw.status_1398.qe;
  assign rcache_line[5][118].status_reg.re    = reg2hw.status_1398.re;


  assign rcache_line[5][119].tag_reg.tag      = reg2hw.tag_1399.q;
  assign rcache_line[5][119].tag_reg.qe       = reg2hw.tag_1399.qe;
  assign rcache_line[5][119].tag_reg.re       = reg2hw.tag_1399.re;
  assign rcache_line[5][119].status_reg.status = reg2hw.status_1399.q;//status_reg_t'(reg2hw.status_1399.q);
  assign rcache_line[5][119].status_reg.qe    = reg2hw.status_1399.qe;
  assign rcache_line[5][119].status_reg.re    = reg2hw.status_1399.re;


  assign rcache_line[5][120].tag_reg.tag      = reg2hw.tag_1400.q;
  assign rcache_line[5][120].tag_reg.qe       = reg2hw.tag_1400.qe;
  assign rcache_line[5][120].tag_reg.re       = reg2hw.tag_1400.re;
  assign rcache_line[5][120].status_reg.status = reg2hw.status_1400.q;//status_reg_t'(reg2hw.status_1400.q);
  assign rcache_line[5][120].status_reg.qe    = reg2hw.status_1400.qe;
  assign rcache_line[5][120].status_reg.re    = reg2hw.status_1400.re;


  assign rcache_line[5][121].tag_reg.tag      = reg2hw.tag_1401.q;
  assign rcache_line[5][121].tag_reg.qe       = reg2hw.tag_1401.qe;
  assign rcache_line[5][121].tag_reg.re       = reg2hw.tag_1401.re;
  assign rcache_line[5][121].status_reg.status = reg2hw.status_1401.q;//status_reg_t'(reg2hw.status_1401.q);
  assign rcache_line[5][121].status_reg.qe    = reg2hw.status_1401.qe;
  assign rcache_line[5][121].status_reg.re    = reg2hw.status_1401.re;


  assign rcache_line[5][122].tag_reg.tag      = reg2hw.tag_1402.q;
  assign rcache_line[5][122].tag_reg.qe       = reg2hw.tag_1402.qe;
  assign rcache_line[5][122].tag_reg.re       = reg2hw.tag_1402.re;
  assign rcache_line[5][122].status_reg.status = reg2hw.status_1402.q;//status_reg_t'(reg2hw.status_1402.q);
  assign rcache_line[5][122].status_reg.qe    = reg2hw.status_1402.qe;
  assign rcache_line[5][122].status_reg.re    = reg2hw.status_1402.re;


  assign rcache_line[5][123].tag_reg.tag      = reg2hw.tag_1403.q;
  assign rcache_line[5][123].tag_reg.qe       = reg2hw.tag_1403.qe;
  assign rcache_line[5][123].tag_reg.re       = reg2hw.tag_1403.re;
  assign rcache_line[5][123].status_reg.status = reg2hw.status_1403.q;//status_reg_t'(reg2hw.status_1403.q);
  assign rcache_line[5][123].status_reg.qe    = reg2hw.status_1403.qe;
  assign rcache_line[5][123].status_reg.re    = reg2hw.status_1403.re;


  assign rcache_line[5][124].tag_reg.tag      = reg2hw.tag_1404.q;
  assign rcache_line[5][124].tag_reg.qe       = reg2hw.tag_1404.qe;
  assign rcache_line[5][124].tag_reg.re       = reg2hw.tag_1404.re;
  assign rcache_line[5][124].status_reg.status = reg2hw.status_1404.q;//status_reg_t'(reg2hw.status_1404.q);
  assign rcache_line[5][124].status_reg.qe    = reg2hw.status_1404.qe;
  assign rcache_line[5][124].status_reg.re    = reg2hw.status_1404.re;


  assign rcache_line[5][125].tag_reg.tag      = reg2hw.tag_1405.q;
  assign rcache_line[5][125].tag_reg.qe       = reg2hw.tag_1405.qe;
  assign rcache_line[5][125].tag_reg.re       = reg2hw.tag_1405.re;
  assign rcache_line[5][125].status_reg.status = reg2hw.status_1405.q;//status_reg_t'(reg2hw.status_1405.q);
  assign rcache_line[5][125].status_reg.qe    = reg2hw.status_1405.qe;
  assign rcache_line[5][125].status_reg.re    = reg2hw.status_1405.re;


  assign rcache_line[5][126].tag_reg.tag      = reg2hw.tag_1406.q;
  assign rcache_line[5][126].tag_reg.qe       = reg2hw.tag_1406.qe;
  assign rcache_line[5][126].tag_reg.re       = reg2hw.tag_1406.re;
  assign rcache_line[5][126].status_reg.status = reg2hw.status_1406.q;//status_reg_t'(reg2hw.status_1406.q);
  assign rcache_line[5][126].status_reg.qe    = reg2hw.status_1406.qe;
  assign rcache_line[5][126].status_reg.re    = reg2hw.status_1406.re;


  assign rcache_line[5][127].tag_reg.tag      = reg2hw.tag_1407.q;
  assign rcache_line[5][127].tag_reg.qe       = reg2hw.tag_1407.qe;
  assign rcache_line[5][127].tag_reg.re       = reg2hw.tag_1407.re;
  assign rcache_line[5][127].status_reg.status = reg2hw.status_1407.q;//status_reg_t'(reg2hw.status_1407.q);
  assign rcache_line[5][127].status_reg.qe    = reg2hw.status_1407.qe;
  assign rcache_line[5][127].status_reg.re    = reg2hw.status_1407.re;


  assign rcache_line[5][128].tag_reg.tag      = reg2hw.tag_1408.q;
  assign rcache_line[5][128].tag_reg.qe       = reg2hw.tag_1408.qe;
  assign rcache_line[5][128].tag_reg.re       = reg2hw.tag_1408.re;
  assign rcache_line[5][128].status_reg.status = reg2hw.status_1408.q;//status_reg_t'(reg2hw.status_1408.q);
  assign rcache_line[5][128].status_reg.qe    = reg2hw.status_1408.qe;
  assign rcache_line[5][128].status_reg.re    = reg2hw.status_1408.re;


  assign rcache_line[5][129].tag_reg.tag      = reg2hw.tag_1409.q;
  assign rcache_line[5][129].tag_reg.qe       = reg2hw.tag_1409.qe;
  assign rcache_line[5][129].tag_reg.re       = reg2hw.tag_1409.re;
  assign rcache_line[5][129].status_reg.status = reg2hw.status_1409.q;//status_reg_t'(reg2hw.status_1409.q);
  assign rcache_line[5][129].status_reg.qe    = reg2hw.status_1409.qe;
  assign rcache_line[5][129].status_reg.re    = reg2hw.status_1409.re;


  assign rcache_line[5][130].tag_reg.tag      = reg2hw.tag_1410.q;
  assign rcache_line[5][130].tag_reg.qe       = reg2hw.tag_1410.qe;
  assign rcache_line[5][130].tag_reg.re       = reg2hw.tag_1410.re;
  assign rcache_line[5][130].status_reg.status = reg2hw.status_1410.q;//status_reg_t'(reg2hw.status_1410.q);
  assign rcache_line[5][130].status_reg.qe    = reg2hw.status_1410.qe;
  assign rcache_line[5][130].status_reg.re    = reg2hw.status_1410.re;


  assign rcache_line[5][131].tag_reg.tag      = reg2hw.tag_1411.q;
  assign rcache_line[5][131].tag_reg.qe       = reg2hw.tag_1411.qe;
  assign rcache_line[5][131].tag_reg.re       = reg2hw.tag_1411.re;
  assign rcache_line[5][131].status_reg.status = reg2hw.status_1411.q;//status_reg_t'(reg2hw.status_1411.q);
  assign rcache_line[5][131].status_reg.qe    = reg2hw.status_1411.qe;
  assign rcache_line[5][131].status_reg.re    = reg2hw.status_1411.re;


  assign rcache_line[5][132].tag_reg.tag      = reg2hw.tag_1412.q;
  assign rcache_line[5][132].tag_reg.qe       = reg2hw.tag_1412.qe;
  assign rcache_line[5][132].tag_reg.re       = reg2hw.tag_1412.re;
  assign rcache_line[5][132].status_reg.status = reg2hw.status_1412.q;//status_reg_t'(reg2hw.status_1412.q);
  assign rcache_line[5][132].status_reg.qe    = reg2hw.status_1412.qe;
  assign rcache_line[5][132].status_reg.re    = reg2hw.status_1412.re;


  assign rcache_line[5][133].tag_reg.tag      = reg2hw.tag_1413.q;
  assign rcache_line[5][133].tag_reg.qe       = reg2hw.tag_1413.qe;
  assign rcache_line[5][133].tag_reg.re       = reg2hw.tag_1413.re;
  assign rcache_line[5][133].status_reg.status = reg2hw.status_1413.q;//status_reg_t'(reg2hw.status_1413.q);
  assign rcache_line[5][133].status_reg.qe    = reg2hw.status_1413.qe;
  assign rcache_line[5][133].status_reg.re    = reg2hw.status_1413.re;


  assign rcache_line[5][134].tag_reg.tag      = reg2hw.tag_1414.q;
  assign rcache_line[5][134].tag_reg.qe       = reg2hw.tag_1414.qe;
  assign rcache_line[5][134].tag_reg.re       = reg2hw.tag_1414.re;
  assign rcache_line[5][134].status_reg.status = reg2hw.status_1414.q;//status_reg_t'(reg2hw.status_1414.q);
  assign rcache_line[5][134].status_reg.qe    = reg2hw.status_1414.qe;
  assign rcache_line[5][134].status_reg.re    = reg2hw.status_1414.re;


  assign rcache_line[5][135].tag_reg.tag      = reg2hw.tag_1415.q;
  assign rcache_line[5][135].tag_reg.qe       = reg2hw.tag_1415.qe;
  assign rcache_line[5][135].tag_reg.re       = reg2hw.tag_1415.re;
  assign rcache_line[5][135].status_reg.status = reg2hw.status_1415.q;//status_reg_t'(reg2hw.status_1415.q);
  assign rcache_line[5][135].status_reg.qe    = reg2hw.status_1415.qe;
  assign rcache_line[5][135].status_reg.re    = reg2hw.status_1415.re;


  assign rcache_line[5][136].tag_reg.tag      = reg2hw.tag_1416.q;
  assign rcache_line[5][136].tag_reg.qe       = reg2hw.tag_1416.qe;
  assign rcache_line[5][136].tag_reg.re       = reg2hw.tag_1416.re;
  assign rcache_line[5][136].status_reg.status = reg2hw.status_1416.q;//status_reg_t'(reg2hw.status_1416.q);
  assign rcache_line[5][136].status_reg.qe    = reg2hw.status_1416.qe;
  assign rcache_line[5][136].status_reg.re    = reg2hw.status_1416.re;


  assign rcache_line[5][137].tag_reg.tag      = reg2hw.tag_1417.q;
  assign rcache_line[5][137].tag_reg.qe       = reg2hw.tag_1417.qe;
  assign rcache_line[5][137].tag_reg.re       = reg2hw.tag_1417.re;
  assign rcache_line[5][137].status_reg.status = reg2hw.status_1417.q;//status_reg_t'(reg2hw.status_1417.q);
  assign rcache_line[5][137].status_reg.qe    = reg2hw.status_1417.qe;
  assign rcache_line[5][137].status_reg.re    = reg2hw.status_1417.re;


  assign rcache_line[5][138].tag_reg.tag      = reg2hw.tag_1418.q;
  assign rcache_line[5][138].tag_reg.qe       = reg2hw.tag_1418.qe;
  assign rcache_line[5][138].tag_reg.re       = reg2hw.tag_1418.re;
  assign rcache_line[5][138].status_reg.status = reg2hw.status_1418.q;//status_reg_t'(reg2hw.status_1418.q);
  assign rcache_line[5][138].status_reg.qe    = reg2hw.status_1418.qe;
  assign rcache_line[5][138].status_reg.re    = reg2hw.status_1418.re;


  assign rcache_line[5][139].tag_reg.tag      = reg2hw.tag_1419.q;
  assign rcache_line[5][139].tag_reg.qe       = reg2hw.tag_1419.qe;
  assign rcache_line[5][139].tag_reg.re       = reg2hw.tag_1419.re;
  assign rcache_line[5][139].status_reg.status = reg2hw.status_1419.q;//status_reg_t'(reg2hw.status_1419.q);
  assign rcache_line[5][139].status_reg.qe    = reg2hw.status_1419.qe;
  assign rcache_line[5][139].status_reg.re    = reg2hw.status_1419.re;


  assign rcache_line[5][140].tag_reg.tag      = reg2hw.tag_1420.q;
  assign rcache_line[5][140].tag_reg.qe       = reg2hw.tag_1420.qe;
  assign rcache_line[5][140].tag_reg.re       = reg2hw.tag_1420.re;
  assign rcache_line[5][140].status_reg.status = reg2hw.status_1420.q;//status_reg_t'(reg2hw.status_1420.q);
  assign rcache_line[5][140].status_reg.qe    = reg2hw.status_1420.qe;
  assign rcache_line[5][140].status_reg.re    = reg2hw.status_1420.re;


  assign rcache_line[5][141].tag_reg.tag      = reg2hw.tag_1421.q;
  assign rcache_line[5][141].tag_reg.qe       = reg2hw.tag_1421.qe;
  assign rcache_line[5][141].tag_reg.re       = reg2hw.tag_1421.re;
  assign rcache_line[5][141].status_reg.status = reg2hw.status_1421.q;//status_reg_t'(reg2hw.status_1421.q);
  assign rcache_line[5][141].status_reg.qe    = reg2hw.status_1421.qe;
  assign rcache_line[5][141].status_reg.re    = reg2hw.status_1421.re;


  assign rcache_line[5][142].tag_reg.tag      = reg2hw.tag_1422.q;
  assign rcache_line[5][142].tag_reg.qe       = reg2hw.tag_1422.qe;
  assign rcache_line[5][142].tag_reg.re       = reg2hw.tag_1422.re;
  assign rcache_line[5][142].status_reg.status = reg2hw.status_1422.q;//status_reg_t'(reg2hw.status_1422.q);
  assign rcache_line[5][142].status_reg.qe    = reg2hw.status_1422.qe;
  assign rcache_line[5][142].status_reg.re    = reg2hw.status_1422.re;


  assign rcache_line[5][143].tag_reg.tag      = reg2hw.tag_1423.q;
  assign rcache_line[5][143].tag_reg.qe       = reg2hw.tag_1423.qe;
  assign rcache_line[5][143].tag_reg.re       = reg2hw.tag_1423.re;
  assign rcache_line[5][143].status_reg.status = reg2hw.status_1423.q;//status_reg_t'(reg2hw.status_1423.q);
  assign rcache_line[5][143].status_reg.qe    = reg2hw.status_1423.qe;
  assign rcache_line[5][143].status_reg.re    = reg2hw.status_1423.re;


  assign rcache_line[5][144].tag_reg.tag      = reg2hw.tag_1424.q;
  assign rcache_line[5][144].tag_reg.qe       = reg2hw.tag_1424.qe;
  assign rcache_line[5][144].tag_reg.re       = reg2hw.tag_1424.re;
  assign rcache_line[5][144].status_reg.status = reg2hw.status_1424.q;//status_reg_t'(reg2hw.status_1424.q);
  assign rcache_line[5][144].status_reg.qe    = reg2hw.status_1424.qe;
  assign rcache_line[5][144].status_reg.re    = reg2hw.status_1424.re;


  assign rcache_line[5][145].tag_reg.tag      = reg2hw.tag_1425.q;
  assign rcache_line[5][145].tag_reg.qe       = reg2hw.tag_1425.qe;
  assign rcache_line[5][145].tag_reg.re       = reg2hw.tag_1425.re;
  assign rcache_line[5][145].status_reg.status = reg2hw.status_1425.q;//status_reg_t'(reg2hw.status_1425.q);
  assign rcache_line[5][145].status_reg.qe    = reg2hw.status_1425.qe;
  assign rcache_line[5][145].status_reg.re    = reg2hw.status_1425.re;


  assign rcache_line[5][146].tag_reg.tag      = reg2hw.tag_1426.q;
  assign rcache_line[5][146].tag_reg.qe       = reg2hw.tag_1426.qe;
  assign rcache_line[5][146].tag_reg.re       = reg2hw.tag_1426.re;
  assign rcache_line[5][146].status_reg.status = reg2hw.status_1426.q;//status_reg_t'(reg2hw.status_1426.q);
  assign rcache_line[5][146].status_reg.qe    = reg2hw.status_1426.qe;
  assign rcache_line[5][146].status_reg.re    = reg2hw.status_1426.re;


  assign rcache_line[5][147].tag_reg.tag      = reg2hw.tag_1427.q;
  assign rcache_line[5][147].tag_reg.qe       = reg2hw.tag_1427.qe;
  assign rcache_line[5][147].tag_reg.re       = reg2hw.tag_1427.re;
  assign rcache_line[5][147].status_reg.status = reg2hw.status_1427.q;//status_reg_t'(reg2hw.status_1427.q);
  assign rcache_line[5][147].status_reg.qe    = reg2hw.status_1427.qe;
  assign rcache_line[5][147].status_reg.re    = reg2hw.status_1427.re;


  assign rcache_line[5][148].tag_reg.tag      = reg2hw.tag_1428.q;
  assign rcache_line[5][148].tag_reg.qe       = reg2hw.tag_1428.qe;
  assign rcache_line[5][148].tag_reg.re       = reg2hw.tag_1428.re;
  assign rcache_line[5][148].status_reg.status = reg2hw.status_1428.q;//status_reg_t'(reg2hw.status_1428.q);
  assign rcache_line[5][148].status_reg.qe    = reg2hw.status_1428.qe;
  assign rcache_line[5][148].status_reg.re    = reg2hw.status_1428.re;


  assign rcache_line[5][149].tag_reg.tag      = reg2hw.tag_1429.q;
  assign rcache_line[5][149].tag_reg.qe       = reg2hw.tag_1429.qe;
  assign rcache_line[5][149].tag_reg.re       = reg2hw.tag_1429.re;
  assign rcache_line[5][149].status_reg.status = reg2hw.status_1429.q;//status_reg_t'(reg2hw.status_1429.q);
  assign rcache_line[5][149].status_reg.qe    = reg2hw.status_1429.qe;
  assign rcache_line[5][149].status_reg.re    = reg2hw.status_1429.re;


  assign rcache_line[5][150].tag_reg.tag      = reg2hw.tag_1430.q;
  assign rcache_line[5][150].tag_reg.qe       = reg2hw.tag_1430.qe;
  assign rcache_line[5][150].tag_reg.re       = reg2hw.tag_1430.re;
  assign rcache_line[5][150].status_reg.status = reg2hw.status_1430.q;//status_reg_t'(reg2hw.status_1430.q);
  assign rcache_line[5][150].status_reg.qe    = reg2hw.status_1430.qe;
  assign rcache_line[5][150].status_reg.re    = reg2hw.status_1430.re;


  assign rcache_line[5][151].tag_reg.tag      = reg2hw.tag_1431.q;
  assign rcache_line[5][151].tag_reg.qe       = reg2hw.tag_1431.qe;
  assign rcache_line[5][151].tag_reg.re       = reg2hw.tag_1431.re;
  assign rcache_line[5][151].status_reg.status = reg2hw.status_1431.q;//status_reg_t'(reg2hw.status_1431.q);
  assign rcache_line[5][151].status_reg.qe    = reg2hw.status_1431.qe;
  assign rcache_line[5][151].status_reg.re    = reg2hw.status_1431.re;


  assign rcache_line[5][152].tag_reg.tag      = reg2hw.tag_1432.q;
  assign rcache_line[5][152].tag_reg.qe       = reg2hw.tag_1432.qe;
  assign rcache_line[5][152].tag_reg.re       = reg2hw.tag_1432.re;
  assign rcache_line[5][152].status_reg.status = reg2hw.status_1432.q;//status_reg_t'(reg2hw.status_1432.q);
  assign rcache_line[5][152].status_reg.qe    = reg2hw.status_1432.qe;
  assign rcache_line[5][152].status_reg.re    = reg2hw.status_1432.re;


  assign rcache_line[5][153].tag_reg.tag      = reg2hw.tag_1433.q;
  assign rcache_line[5][153].tag_reg.qe       = reg2hw.tag_1433.qe;
  assign rcache_line[5][153].tag_reg.re       = reg2hw.tag_1433.re;
  assign rcache_line[5][153].status_reg.status = reg2hw.status_1433.q;//status_reg_t'(reg2hw.status_1433.q);
  assign rcache_line[5][153].status_reg.qe    = reg2hw.status_1433.qe;
  assign rcache_line[5][153].status_reg.re    = reg2hw.status_1433.re;


  assign rcache_line[5][154].tag_reg.tag      = reg2hw.tag_1434.q;
  assign rcache_line[5][154].tag_reg.qe       = reg2hw.tag_1434.qe;
  assign rcache_line[5][154].tag_reg.re       = reg2hw.tag_1434.re;
  assign rcache_line[5][154].status_reg.status = reg2hw.status_1434.q;//status_reg_t'(reg2hw.status_1434.q);
  assign rcache_line[5][154].status_reg.qe    = reg2hw.status_1434.qe;
  assign rcache_line[5][154].status_reg.re    = reg2hw.status_1434.re;


  assign rcache_line[5][155].tag_reg.tag      = reg2hw.tag_1435.q;
  assign rcache_line[5][155].tag_reg.qe       = reg2hw.tag_1435.qe;
  assign rcache_line[5][155].tag_reg.re       = reg2hw.tag_1435.re;
  assign rcache_line[5][155].status_reg.status = reg2hw.status_1435.q;//status_reg_t'(reg2hw.status_1435.q);
  assign rcache_line[5][155].status_reg.qe    = reg2hw.status_1435.qe;
  assign rcache_line[5][155].status_reg.re    = reg2hw.status_1435.re;


  assign rcache_line[5][156].tag_reg.tag      = reg2hw.tag_1436.q;
  assign rcache_line[5][156].tag_reg.qe       = reg2hw.tag_1436.qe;
  assign rcache_line[5][156].tag_reg.re       = reg2hw.tag_1436.re;
  assign rcache_line[5][156].status_reg.status = reg2hw.status_1436.q;//status_reg_t'(reg2hw.status_1436.q);
  assign rcache_line[5][156].status_reg.qe    = reg2hw.status_1436.qe;
  assign rcache_line[5][156].status_reg.re    = reg2hw.status_1436.re;


  assign rcache_line[5][157].tag_reg.tag      = reg2hw.tag_1437.q;
  assign rcache_line[5][157].tag_reg.qe       = reg2hw.tag_1437.qe;
  assign rcache_line[5][157].tag_reg.re       = reg2hw.tag_1437.re;
  assign rcache_line[5][157].status_reg.status = reg2hw.status_1437.q;//status_reg_t'(reg2hw.status_1437.q);
  assign rcache_line[5][157].status_reg.qe    = reg2hw.status_1437.qe;
  assign rcache_line[5][157].status_reg.re    = reg2hw.status_1437.re;


  assign rcache_line[5][158].tag_reg.tag      = reg2hw.tag_1438.q;
  assign rcache_line[5][158].tag_reg.qe       = reg2hw.tag_1438.qe;
  assign rcache_line[5][158].tag_reg.re       = reg2hw.tag_1438.re;
  assign rcache_line[5][158].status_reg.status = reg2hw.status_1438.q;//status_reg_t'(reg2hw.status_1438.q);
  assign rcache_line[5][158].status_reg.qe    = reg2hw.status_1438.qe;
  assign rcache_line[5][158].status_reg.re    = reg2hw.status_1438.re;


  assign rcache_line[5][159].tag_reg.tag      = reg2hw.tag_1439.q;
  assign rcache_line[5][159].tag_reg.qe       = reg2hw.tag_1439.qe;
  assign rcache_line[5][159].tag_reg.re       = reg2hw.tag_1439.re;
  assign rcache_line[5][159].status_reg.status = reg2hw.status_1439.q;//status_reg_t'(reg2hw.status_1439.q);
  assign rcache_line[5][159].status_reg.qe    = reg2hw.status_1439.qe;
  assign rcache_line[5][159].status_reg.re    = reg2hw.status_1439.re;


  assign rcache_line[5][160].tag_reg.tag      = reg2hw.tag_1440.q;
  assign rcache_line[5][160].tag_reg.qe       = reg2hw.tag_1440.qe;
  assign rcache_line[5][160].tag_reg.re       = reg2hw.tag_1440.re;
  assign rcache_line[5][160].status_reg.status = reg2hw.status_1440.q;//status_reg_t'(reg2hw.status_1440.q);
  assign rcache_line[5][160].status_reg.qe    = reg2hw.status_1440.qe;
  assign rcache_line[5][160].status_reg.re    = reg2hw.status_1440.re;


  assign rcache_line[5][161].tag_reg.tag      = reg2hw.tag_1441.q;
  assign rcache_line[5][161].tag_reg.qe       = reg2hw.tag_1441.qe;
  assign rcache_line[5][161].tag_reg.re       = reg2hw.tag_1441.re;
  assign rcache_line[5][161].status_reg.status = reg2hw.status_1441.q;//status_reg_t'(reg2hw.status_1441.q);
  assign rcache_line[5][161].status_reg.qe    = reg2hw.status_1441.qe;
  assign rcache_line[5][161].status_reg.re    = reg2hw.status_1441.re;


  assign rcache_line[5][162].tag_reg.tag      = reg2hw.tag_1442.q;
  assign rcache_line[5][162].tag_reg.qe       = reg2hw.tag_1442.qe;
  assign rcache_line[5][162].tag_reg.re       = reg2hw.tag_1442.re;
  assign rcache_line[5][162].status_reg.status = reg2hw.status_1442.q;//status_reg_t'(reg2hw.status_1442.q);
  assign rcache_line[5][162].status_reg.qe    = reg2hw.status_1442.qe;
  assign rcache_line[5][162].status_reg.re    = reg2hw.status_1442.re;


  assign rcache_line[5][163].tag_reg.tag      = reg2hw.tag_1443.q;
  assign rcache_line[5][163].tag_reg.qe       = reg2hw.tag_1443.qe;
  assign rcache_line[5][163].tag_reg.re       = reg2hw.tag_1443.re;
  assign rcache_line[5][163].status_reg.status = reg2hw.status_1443.q;//status_reg_t'(reg2hw.status_1443.q);
  assign rcache_line[5][163].status_reg.qe    = reg2hw.status_1443.qe;
  assign rcache_line[5][163].status_reg.re    = reg2hw.status_1443.re;


  assign rcache_line[5][164].tag_reg.tag      = reg2hw.tag_1444.q;
  assign rcache_line[5][164].tag_reg.qe       = reg2hw.tag_1444.qe;
  assign rcache_line[5][164].tag_reg.re       = reg2hw.tag_1444.re;
  assign rcache_line[5][164].status_reg.status = reg2hw.status_1444.q;//status_reg_t'(reg2hw.status_1444.q);
  assign rcache_line[5][164].status_reg.qe    = reg2hw.status_1444.qe;
  assign rcache_line[5][164].status_reg.re    = reg2hw.status_1444.re;


  assign rcache_line[5][165].tag_reg.tag      = reg2hw.tag_1445.q;
  assign rcache_line[5][165].tag_reg.qe       = reg2hw.tag_1445.qe;
  assign rcache_line[5][165].tag_reg.re       = reg2hw.tag_1445.re;
  assign rcache_line[5][165].status_reg.status = reg2hw.status_1445.q;//status_reg_t'(reg2hw.status_1445.q);
  assign rcache_line[5][165].status_reg.qe    = reg2hw.status_1445.qe;
  assign rcache_line[5][165].status_reg.re    = reg2hw.status_1445.re;


  assign rcache_line[5][166].tag_reg.tag      = reg2hw.tag_1446.q;
  assign rcache_line[5][166].tag_reg.qe       = reg2hw.tag_1446.qe;
  assign rcache_line[5][166].tag_reg.re       = reg2hw.tag_1446.re;
  assign rcache_line[5][166].status_reg.status = reg2hw.status_1446.q;//status_reg_t'(reg2hw.status_1446.q);
  assign rcache_line[5][166].status_reg.qe    = reg2hw.status_1446.qe;
  assign rcache_line[5][166].status_reg.re    = reg2hw.status_1446.re;


  assign rcache_line[5][167].tag_reg.tag      = reg2hw.tag_1447.q;
  assign rcache_line[5][167].tag_reg.qe       = reg2hw.tag_1447.qe;
  assign rcache_line[5][167].tag_reg.re       = reg2hw.tag_1447.re;
  assign rcache_line[5][167].status_reg.status = reg2hw.status_1447.q;//status_reg_t'(reg2hw.status_1447.q);
  assign rcache_line[5][167].status_reg.qe    = reg2hw.status_1447.qe;
  assign rcache_line[5][167].status_reg.re    = reg2hw.status_1447.re;


  assign rcache_line[5][168].tag_reg.tag      = reg2hw.tag_1448.q;
  assign rcache_line[5][168].tag_reg.qe       = reg2hw.tag_1448.qe;
  assign rcache_line[5][168].tag_reg.re       = reg2hw.tag_1448.re;
  assign rcache_line[5][168].status_reg.status = reg2hw.status_1448.q;//status_reg_t'(reg2hw.status_1448.q);
  assign rcache_line[5][168].status_reg.qe    = reg2hw.status_1448.qe;
  assign rcache_line[5][168].status_reg.re    = reg2hw.status_1448.re;


  assign rcache_line[5][169].tag_reg.tag      = reg2hw.tag_1449.q;
  assign rcache_line[5][169].tag_reg.qe       = reg2hw.tag_1449.qe;
  assign rcache_line[5][169].tag_reg.re       = reg2hw.tag_1449.re;
  assign rcache_line[5][169].status_reg.status = reg2hw.status_1449.q;//status_reg_t'(reg2hw.status_1449.q);
  assign rcache_line[5][169].status_reg.qe    = reg2hw.status_1449.qe;
  assign rcache_line[5][169].status_reg.re    = reg2hw.status_1449.re;


  assign rcache_line[5][170].tag_reg.tag      = reg2hw.tag_1450.q;
  assign rcache_line[5][170].tag_reg.qe       = reg2hw.tag_1450.qe;
  assign rcache_line[5][170].tag_reg.re       = reg2hw.tag_1450.re;
  assign rcache_line[5][170].status_reg.status = reg2hw.status_1450.q;//status_reg_t'(reg2hw.status_1450.q);
  assign rcache_line[5][170].status_reg.qe    = reg2hw.status_1450.qe;
  assign rcache_line[5][170].status_reg.re    = reg2hw.status_1450.re;


  assign rcache_line[5][171].tag_reg.tag      = reg2hw.tag_1451.q;
  assign rcache_line[5][171].tag_reg.qe       = reg2hw.tag_1451.qe;
  assign rcache_line[5][171].tag_reg.re       = reg2hw.tag_1451.re;
  assign rcache_line[5][171].status_reg.status = reg2hw.status_1451.q;//status_reg_t'(reg2hw.status_1451.q);
  assign rcache_line[5][171].status_reg.qe    = reg2hw.status_1451.qe;
  assign rcache_line[5][171].status_reg.re    = reg2hw.status_1451.re;


  assign rcache_line[5][172].tag_reg.tag      = reg2hw.tag_1452.q;
  assign rcache_line[5][172].tag_reg.qe       = reg2hw.tag_1452.qe;
  assign rcache_line[5][172].tag_reg.re       = reg2hw.tag_1452.re;
  assign rcache_line[5][172].status_reg.status = reg2hw.status_1452.q;//status_reg_t'(reg2hw.status_1452.q);
  assign rcache_line[5][172].status_reg.qe    = reg2hw.status_1452.qe;
  assign rcache_line[5][172].status_reg.re    = reg2hw.status_1452.re;


  assign rcache_line[5][173].tag_reg.tag      = reg2hw.tag_1453.q;
  assign rcache_line[5][173].tag_reg.qe       = reg2hw.tag_1453.qe;
  assign rcache_line[5][173].tag_reg.re       = reg2hw.tag_1453.re;
  assign rcache_line[5][173].status_reg.status = reg2hw.status_1453.q;//status_reg_t'(reg2hw.status_1453.q);
  assign rcache_line[5][173].status_reg.qe    = reg2hw.status_1453.qe;
  assign rcache_line[5][173].status_reg.re    = reg2hw.status_1453.re;


  assign rcache_line[5][174].tag_reg.tag      = reg2hw.tag_1454.q;
  assign rcache_line[5][174].tag_reg.qe       = reg2hw.tag_1454.qe;
  assign rcache_line[5][174].tag_reg.re       = reg2hw.tag_1454.re;
  assign rcache_line[5][174].status_reg.status = reg2hw.status_1454.q;//status_reg_t'(reg2hw.status_1454.q);
  assign rcache_line[5][174].status_reg.qe    = reg2hw.status_1454.qe;
  assign rcache_line[5][174].status_reg.re    = reg2hw.status_1454.re;


  assign rcache_line[5][175].tag_reg.tag      = reg2hw.tag_1455.q;
  assign rcache_line[5][175].tag_reg.qe       = reg2hw.tag_1455.qe;
  assign rcache_line[5][175].tag_reg.re       = reg2hw.tag_1455.re;
  assign rcache_line[5][175].status_reg.status = reg2hw.status_1455.q;//status_reg_t'(reg2hw.status_1455.q);
  assign rcache_line[5][175].status_reg.qe    = reg2hw.status_1455.qe;
  assign rcache_line[5][175].status_reg.re    = reg2hw.status_1455.re;


  assign rcache_line[5][176].tag_reg.tag      = reg2hw.tag_1456.q;
  assign rcache_line[5][176].tag_reg.qe       = reg2hw.tag_1456.qe;
  assign rcache_line[5][176].tag_reg.re       = reg2hw.tag_1456.re;
  assign rcache_line[5][176].status_reg.status = reg2hw.status_1456.q;//status_reg_t'(reg2hw.status_1456.q);
  assign rcache_line[5][176].status_reg.qe    = reg2hw.status_1456.qe;
  assign rcache_line[5][176].status_reg.re    = reg2hw.status_1456.re;


  assign rcache_line[5][177].tag_reg.tag      = reg2hw.tag_1457.q;
  assign rcache_line[5][177].tag_reg.qe       = reg2hw.tag_1457.qe;
  assign rcache_line[5][177].tag_reg.re       = reg2hw.tag_1457.re;
  assign rcache_line[5][177].status_reg.status = reg2hw.status_1457.q;//status_reg_t'(reg2hw.status_1457.q);
  assign rcache_line[5][177].status_reg.qe    = reg2hw.status_1457.qe;
  assign rcache_line[5][177].status_reg.re    = reg2hw.status_1457.re;


  assign rcache_line[5][178].tag_reg.tag      = reg2hw.tag_1458.q;
  assign rcache_line[5][178].tag_reg.qe       = reg2hw.tag_1458.qe;
  assign rcache_line[5][178].tag_reg.re       = reg2hw.tag_1458.re;
  assign rcache_line[5][178].status_reg.status = reg2hw.status_1458.q;//status_reg_t'(reg2hw.status_1458.q);
  assign rcache_line[5][178].status_reg.qe    = reg2hw.status_1458.qe;
  assign rcache_line[5][178].status_reg.re    = reg2hw.status_1458.re;


  assign rcache_line[5][179].tag_reg.tag      = reg2hw.tag_1459.q;
  assign rcache_line[5][179].tag_reg.qe       = reg2hw.tag_1459.qe;
  assign rcache_line[5][179].tag_reg.re       = reg2hw.tag_1459.re;
  assign rcache_line[5][179].status_reg.status = reg2hw.status_1459.q;//status_reg_t'(reg2hw.status_1459.q);
  assign rcache_line[5][179].status_reg.qe    = reg2hw.status_1459.qe;
  assign rcache_line[5][179].status_reg.re    = reg2hw.status_1459.re;


  assign rcache_line[5][180].tag_reg.tag      = reg2hw.tag_1460.q;
  assign rcache_line[5][180].tag_reg.qe       = reg2hw.tag_1460.qe;
  assign rcache_line[5][180].tag_reg.re       = reg2hw.tag_1460.re;
  assign rcache_line[5][180].status_reg.status = reg2hw.status_1460.q;//status_reg_t'(reg2hw.status_1460.q);
  assign rcache_line[5][180].status_reg.qe    = reg2hw.status_1460.qe;
  assign rcache_line[5][180].status_reg.re    = reg2hw.status_1460.re;


  assign rcache_line[5][181].tag_reg.tag      = reg2hw.tag_1461.q;
  assign rcache_line[5][181].tag_reg.qe       = reg2hw.tag_1461.qe;
  assign rcache_line[5][181].tag_reg.re       = reg2hw.tag_1461.re;
  assign rcache_line[5][181].status_reg.status = reg2hw.status_1461.q;//status_reg_t'(reg2hw.status_1461.q);
  assign rcache_line[5][181].status_reg.qe    = reg2hw.status_1461.qe;
  assign rcache_line[5][181].status_reg.re    = reg2hw.status_1461.re;


  assign rcache_line[5][182].tag_reg.tag      = reg2hw.tag_1462.q;
  assign rcache_line[5][182].tag_reg.qe       = reg2hw.tag_1462.qe;
  assign rcache_line[5][182].tag_reg.re       = reg2hw.tag_1462.re;
  assign rcache_line[5][182].status_reg.status = reg2hw.status_1462.q;//status_reg_t'(reg2hw.status_1462.q);
  assign rcache_line[5][182].status_reg.qe    = reg2hw.status_1462.qe;
  assign rcache_line[5][182].status_reg.re    = reg2hw.status_1462.re;


  assign rcache_line[5][183].tag_reg.tag      = reg2hw.tag_1463.q;
  assign rcache_line[5][183].tag_reg.qe       = reg2hw.tag_1463.qe;
  assign rcache_line[5][183].tag_reg.re       = reg2hw.tag_1463.re;
  assign rcache_line[5][183].status_reg.status = reg2hw.status_1463.q;//status_reg_t'(reg2hw.status_1463.q);
  assign rcache_line[5][183].status_reg.qe    = reg2hw.status_1463.qe;
  assign rcache_line[5][183].status_reg.re    = reg2hw.status_1463.re;


  assign rcache_line[5][184].tag_reg.tag      = reg2hw.tag_1464.q;
  assign rcache_line[5][184].tag_reg.qe       = reg2hw.tag_1464.qe;
  assign rcache_line[5][184].tag_reg.re       = reg2hw.tag_1464.re;
  assign rcache_line[5][184].status_reg.status = reg2hw.status_1464.q;//status_reg_t'(reg2hw.status_1464.q);
  assign rcache_line[5][184].status_reg.qe    = reg2hw.status_1464.qe;
  assign rcache_line[5][184].status_reg.re    = reg2hw.status_1464.re;


  assign rcache_line[5][185].tag_reg.tag      = reg2hw.tag_1465.q;
  assign rcache_line[5][185].tag_reg.qe       = reg2hw.tag_1465.qe;
  assign rcache_line[5][185].tag_reg.re       = reg2hw.tag_1465.re;
  assign rcache_line[5][185].status_reg.status = reg2hw.status_1465.q;//status_reg_t'(reg2hw.status_1465.q);
  assign rcache_line[5][185].status_reg.qe    = reg2hw.status_1465.qe;
  assign rcache_line[5][185].status_reg.re    = reg2hw.status_1465.re;


  assign rcache_line[5][186].tag_reg.tag      = reg2hw.tag_1466.q;
  assign rcache_line[5][186].tag_reg.qe       = reg2hw.tag_1466.qe;
  assign rcache_line[5][186].tag_reg.re       = reg2hw.tag_1466.re;
  assign rcache_line[5][186].status_reg.status = reg2hw.status_1466.q;//status_reg_t'(reg2hw.status_1466.q);
  assign rcache_line[5][186].status_reg.qe    = reg2hw.status_1466.qe;
  assign rcache_line[5][186].status_reg.re    = reg2hw.status_1466.re;


  assign rcache_line[5][187].tag_reg.tag      = reg2hw.tag_1467.q;
  assign rcache_line[5][187].tag_reg.qe       = reg2hw.tag_1467.qe;
  assign rcache_line[5][187].tag_reg.re       = reg2hw.tag_1467.re;
  assign rcache_line[5][187].status_reg.status = reg2hw.status_1467.q;//status_reg_t'(reg2hw.status_1467.q);
  assign rcache_line[5][187].status_reg.qe    = reg2hw.status_1467.qe;
  assign rcache_line[5][187].status_reg.re    = reg2hw.status_1467.re;


  assign rcache_line[5][188].tag_reg.tag      = reg2hw.tag_1468.q;
  assign rcache_line[5][188].tag_reg.qe       = reg2hw.tag_1468.qe;
  assign rcache_line[5][188].tag_reg.re       = reg2hw.tag_1468.re;
  assign rcache_line[5][188].status_reg.status = reg2hw.status_1468.q;//status_reg_t'(reg2hw.status_1468.q);
  assign rcache_line[5][188].status_reg.qe    = reg2hw.status_1468.qe;
  assign rcache_line[5][188].status_reg.re    = reg2hw.status_1468.re;


  assign rcache_line[5][189].tag_reg.tag      = reg2hw.tag_1469.q;
  assign rcache_line[5][189].tag_reg.qe       = reg2hw.tag_1469.qe;
  assign rcache_line[5][189].tag_reg.re       = reg2hw.tag_1469.re;
  assign rcache_line[5][189].status_reg.status = reg2hw.status_1469.q;//status_reg_t'(reg2hw.status_1469.q);
  assign rcache_line[5][189].status_reg.qe    = reg2hw.status_1469.qe;
  assign rcache_line[5][189].status_reg.re    = reg2hw.status_1469.re;


  assign rcache_line[5][190].tag_reg.tag      = reg2hw.tag_1470.q;
  assign rcache_line[5][190].tag_reg.qe       = reg2hw.tag_1470.qe;
  assign rcache_line[5][190].tag_reg.re       = reg2hw.tag_1470.re;
  assign rcache_line[5][190].status_reg.status = reg2hw.status_1470.q;//status_reg_t'(reg2hw.status_1470.q);
  assign rcache_line[5][190].status_reg.qe    = reg2hw.status_1470.qe;
  assign rcache_line[5][190].status_reg.re    = reg2hw.status_1470.re;


  assign rcache_line[5][191].tag_reg.tag      = reg2hw.tag_1471.q;
  assign rcache_line[5][191].tag_reg.qe       = reg2hw.tag_1471.qe;
  assign rcache_line[5][191].tag_reg.re       = reg2hw.tag_1471.re;
  assign rcache_line[5][191].status_reg.status = reg2hw.status_1471.q;//status_reg_t'(reg2hw.status_1471.q);
  assign rcache_line[5][191].status_reg.qe    = reg2hw.status_1471.qe;
  assign rcache_line[5][191].status_reg.re    = reg2hw.status_1471.re;


  assign rcache_line[5][192].tag_reg.tag      = reg2hw.tag_1472.q;
  assign rcache_line[5][192].tag_reg.qe       = reg2hw.tag_1472.qe;
  assign rcache_line[5][192].tag_reg.re       = reg2hw.tag_1472.re;
  assign rcache_line[5][192].status_reg.status = reg2hw.status_1472.q;//status_reg_t'(reg2hw.status_1472.q);
  assign rcache_line[5][192].status_reg.qe    = reg2hw.status_1472.qe;
  assign rcache_line[5][192].status_reg.re    = reg2hw.status_1472.re;


  assign rcache_line[5][193].tag_reg.tag      = reg2hw.tag_1473.q;
  assign rcache_line[5][193].tag_reg.qe       = reg2hw.tag_1473.qe;
  assign rcache_line[5][193].tag_reg.re       = reg2hw.tag_1473.re;
  assign rcache_line[5][193].status_reg.status = reg2hw.status_1473.q;//status_reg_t'(reg2hw.status_1473.q);
  assign rcache_line[5][193].status_reg.qe    = reg2hw.status_1473.qe;
  assign rcache_line[5][193].status_reg.re    = reg2hw.status_1473.re;


  assign rcache_line[5][194].tag_reg.tag      = reg2hw.tag_1474.q;
  assign rcache_line[5][194].tag_reg.qe       = reg2hw.tag_1474.qe;
  assign rcache_line[5][194].tag_reg.re       = reg2hw.tag_1474.re;
  assign rcache_line[5][194].status_reg.status = reg2hw.status_1474.q;//status_reg_t'(reg2hw.status_1474.q);
  assign rcache_line[5][194].status_reg.qe    = reg2hw.status_1474.qe;
  assign rcache_line[5][194].status_reg.re    = reg2hw.status_1474.re;


  assign rcache_line[5][195].tag_reg.tag      = reg2hw.tag_1475.q;
  assign rcache_line[5][195].tag_reg.qe       = reg2hw.tag_1475.qe;
  assign rcache_line[5][195].tag_reg.re       = reg2hw.tag_1475.re;
  assign rcache_line[5][195].status_reg.status = reg2hw.status_1475.q;//status_reg_t'(reg2hw.status_1475.q);
  assign rcache_line[5][195].status_reg.qe    = reg2hw.status_1475.qe;
  assign rcache_line[5][195].status_reg.re    = reg2hw.status_1475.re;


  assign rcache_line[5][196].tag_reg.tag      = reg2hw.tag_1476.q;
  assign rcache_line[5][196].tag_reg.qe       = reg2hw.tag_1476.qe;
  assign rcache_line[5][196].tag_reg.re       = reg2hw.tag_1476.re;
  assign rcache_line[5][196].status_reg.status = reg2hw.status_1476.q;//status_reg_t'(reg2hw.status_1476.q);
  assign rcache_line[5][196].status_reg.qe    = reg2hw.status_1476.qe;
  assign rcache_line[5][196].status_reg.re    = reg2hw.status_1476.re;


  assign rcache_line[5][197].tag_reg.tag      = reg2hw.tag_1477.q;
  assign rcache_line[5][197].tag_reg.qe       = reg2hw.tag_1477.qe;
  assign rcache_line[5][197].tag_reg.re       = reg2hw.tag_1477.re;
  assign rcache_line[5][197].status_reg.status = reg2hw.status_1477.q;//status_reg_t'(reg2hw.status_1477.q);
  assign rcache_line[5][197].status_reg.qe    = reg2hw.status_1477.qe;
  assign rcache_line[5][197].status_reg.re    = reg2hw.status_1477.re;


  assign rcache_line[5][198].tag_reg.tag      = reg2hw.tag_1478.q;
  assign rcache_line[5][198].tag_reg.qe       = reg2hw.tag_1478.qe;
  assign rcache_line[5][198].tag_reg.re       = reg2hw.tag_1478.re;
  assign rcache_line[5][198].status_reg.status = reg2hw.status_1478.q;//status_reg_t'(reg2hw.status_1478.q);
  assign rcache_line[5][198].status_reg.qe    = reg2hw.status_1478.qe;
  assign rcache_line[5][198].status_reg.re    = reg2hw.status_1478.re;


  assign rcache_line[5][199].tag_reg.tag      = reg2hw.tag_1479.q;
  assign rcache_line[5][199].tag_reg.qe       = reg2hw.tag_1479.qe;
  assign rcache_line[5][199].tag_reg.re       = reg2hw.tag_1479.re;
  assign rcache_line[5][199].status_reg.status = reg2hw.status_1479.q;//status_reg_t'(reg2hw.status_1479.q);
  assign rcache_line[5][199].status_reg.qe    = reg2hw.status_1479.qe;
  assign rcache_line[5][199].status_reg.re    = reg2hw.status_1479.re;


  assign rcache_line[5][200].tag_reg.tag      = reg2hw.tag_1480.q;
  assign rcache_line[5][200].tag_reg.qe       = reg2hw.tag_1480.qe;
  assign rcache_line[5][200].tag_reg.re       = reg2hw.tag_1480.re;
  assign rcache_line[5][200].status_reg.status = reg2hw.status_1480.q;//status_reg_t'(reg2hw.status_1480.q);
  assign rcache_line[5][200].status_reg.qe    = reg2hw.status_1480.qe;
  assign rcache_line[5][200].status_reg.re    = reg2hw.status_1480.re;


  assign rcache_line[5][201].tag_reg.tag      = reg2hw.tag_1481.q;
  assign rcache_line[5][201].tag_reg.qe       = reg2hw.tag_1481.qe;
  assign rcache_line[5][201].tag_reg.re       = reg2hw.tag_1481.re;
  assign rcache_line[5][201].status_reg.status = reg2hw.status_1481.q;//status_reg_t'(reg2hw.status_1481.q);
  assign rcache_line[5][201].status_reg.qe    = reg2hw.status_1481.qe;
  assign rcache_line[5][201].status_reg.re    = reg2hw.status_1481.re;


  assign rcache_line[5][202].tag_reg.tag      = reg2hw.tag_1482.q;
  assign rcache_line[5][202].tag_reg.qe       = reg2hw.tag_1482.qe;
  assign rcache_line[5][202].tag_reg.re       = reg2hw.tag_1482.re;
  assign rcache_line[5][202].status_reg.status = reg2hw.status_1482.q;//status_reg_t'(reg2hw.status_1482.q);
  assign rcache_line[5][202].status_reg.qe    = reg2hw.status_1482.qe;
  assign rcache_line[5][202].status_reg.re    = reg2hw.status_1482.re;


  assign rcache_line[5][203].tag_reg.tag      = reg2hw.tag_1483.q;
  assign rcache_line[5][203].tag_reg.qe       = reg2hw.tag_1483.qe;
  assign rcache_line[5][203].tag_reg.re       = reg2hw.tag_1483.re;
  assign rcache_line[5][203].status_reg.status = reg2hw.status_1483.q;//status_reg_t'(reg2hw.status_1483.q);
  assign rcache_line[5][203].status_reg.qe    = reg2hw.status_1483.qe;
  assign rcache_line[5][203].status_reg.re    = reg2hw.status_1483.re;


  assign rcache_line[5][204].tag_reg.tag      = reg2hw.tag_1484.q;
  assign rcache_line[5][204].tag_reg.qe       = reg2hw.tag_1484.qe;
  assign rcache_line[5][204].tag_reg.re       = reg2hw.tag_1484.re;
  assign rcache_line[5][204].status_reg.status = reg2hw.status_1484.q;//status_reg_t'(reg2hw.status_1484.q);
  assign rcache_line[5][204].status_reg.qe    = reg2hw.status_1484.qe;
  assign rcache_line[5][204].status_reg.re    = reg2hw.status_1484.re;


  assign rcache_line[5][205].tag_reg.tag      = reg2hw.tag_1485.q;
  assign rcache_line[5][205].tag_reg.qe       = reg2hw.tag_1485.qe;
  assign rcache_line[5][205].tag_reg.re       = reg2hw.tag_1485.re;
  assign rcache_line[5][205].status_reg.status = reg2hw.status_1485.q;//status_reg_t'(reg2hw.status_1485.q);
  assign rcache_line[5][205].status_reg.qe    = reg2hw.status_1485.qe;
  assign rcache_line[5][205].status_reg.re    = reg2hw.status_1485.re;


  assign rcache_line[5][206].tag_reg.tag      = reg2hw.tag_1486.q;
  assign rcache_line[5][206].tag_reg.qe       = reg2hw.tag_1486.qe;
  assign rcache_line[5][206].tag_reg.re       = reg2hw.tag_1486.re;
  assign rcache_line[5][206].status_reg.status = reg2hw.status_1486.q;//status_reg_t'(reg2hw.status_1486.q);
  assign rcache_line[5][206].status_reg.qe    = reg2hw.status_1486.qe;
  assign rcache_line[5][206].status_reg.re    = reg2hw.status_1486.re;


  assign rcache_line[5][207].tag_reg.tag      = reg2hw.tag_1487.q;
  assign rcache_line[5][207].tag_reg.qe       = reg2hw.tag_1487.qe;
  assign rcache_line[5][207].tag_reg.re       = reg2hw.tag_1487.re;
  assign rcache_line[5][207].status_reg.status = reg2hw.status_1487.q;//status_reg_t'(reg2hw.status_1487.q);
  assign rcache_line[5][207].status_reg.qe    = reg2hw.status_1487.qe;
  assign rcache_line[5][207].status_reg.re    = reg2hw.status_1487.re;


  assign rcache_line[5][208].tag_reg.tag      = reg2hw.tag_1488.q;
  assign rcache_line[5][208].tag_reg.qe       = reg2hw.tag_1488.qe;
  assign rcache_line[5][208].tag_reg.re       = reg2hw.tag_1488.re;
  assign rcache_line[5][208].status_reg.status = reg2hw.status_1488.q;//status_reg_t'(reg2hw.status_1488.q);
  assign rcache_line[5][208].status_reg.qe    = reg2hw.status_1488.qe;
  assign rcache_line[5][208].status_reg.re    = reg2hw.status_1488.re;


  assign rcache_line[5][209].tag_reg.tag      = reg2hw.tag_1489.q;
  assign rcache_line[5][209].tag_reg.qe       = reg2hw.tag_1489.qe;
  assign rcache_line[5][209].tag_reg.re       = reg2hw.tag_1489.re;
  assign rcache_line[5][209].status_reg.status = reg2hw.status_1489.q;//status_reg_t'(reg2hw.status_1489.q);
  assign rcache_line[5][209].status_reg.qe    = reg2hw.status_1489.qe;
  assign rcache_line[5][209].status_reg.re    = reg2hw.status_1489.re;


  assign rcache_line[5][210].tag_reg.tag      = reg2hw.tag_1490.q;
  assign rcache_line[5][210].tag_reg.qe       = reg2hw.tag_1490.qe;
  assign rcache_line[5][210].tag_reg.re       = reg2hw.tag_1490.re;
  assign rcache_line[5][210].status_reg.status = reg2hw.status_1490.q;//status_reg_t'(reg2hw.status_1490.q);
  assign rcache_line[5][210].status_reg.qe    = reg2hw.status_1490.qe;
  assign rcache_line[5][210].status_reg.re    = reg2hw.status_1490.re;


  assign rcache_line[5][211].tag_reg.tag      = reg2hw.tag_1491.q;
  assign rcache_line[5][211].tag_reg.qe       = reg2hw.tag_1491.qe;
  assign rcache_line[5][211].tag_reg.re       = reg2hw.tag_1491.re;
  assign rcache_line[5][211].status_reg.status = reg2hw.status_1491.q;//status_reg_t'(reg2hw.status_1491.q);
  assign rcache_line[5][211].status_reg.qe    = reg2hw.status_1491.qe;
  assign rcache_line[5][211].status_reg.re    = reg2hw.status_1491.re;


  assign rcache_line[5][212].tag_reg.tag      = reg2hw.tag_1492.q;
  assign rcache_line[5][212].tag_reg.qe       = reg2hw.tag_1492.qe;
  assign rcache_line[5][212].tag_reg.re       = reg2hw.tag_1492.re;
  assign rcache_line[5][212].status_reg.status = reg2hw.status_1492.q;//status_reg_t'(reg2hw.status_1492.q);
  assign rcache_line[5][212].status_reg.qe    = reg2hw.status_1492.qe;
  assign rcache_line[5][212].status_reg.re    = reg2hw.status_1492.re;


  assign rcache_line[5][213].tag_reg.tag      = reg2hw.tag_1493.q;
  assign rcache_line[5][213].tag_reg.qe       = reg2hw.tag_1493.qe;
  assign rcache_line[5][213].tag_reg.re       = reg2hw.tag_1493.re;
  assign rcache_line[5][213].status_reg.status = reg2hw.status_1493.q;//status_reg_t'(reg2hw.status_1493.q);
  assign rcache_line[5][213].status_reg.qe    = reg2hw.status_1493.qe;
  assign rcache_line[5][213].status_reg.re    = reg2hw.status_1493.re;


  assign rcache_line[5][214].tag_reg.tag      = reg2hw.tag_1494.q;
  assign rcache_line[5][214].tag_reg.qe       = reg2hw.tag_1494.qe;
  assign rcache_line[5][214].tag_reg.re       = reg2hw.tag_1494.re;
  assign rcache_line[5][214].status_reg.status = reg2hw.status_1494.q;//status_reg_t'(reg2hw.status_1494.q);
  assign rcache_line[5][214].status_reg.qe    = reg2hw.status_1494.qe;
  assign rcache_line[5][214].status_reg.re    = reg2hw.status_1494.re;


  assign rcache_line[5][215].tag_reg.tag      = reg2hw.tag_1495.q;
  assign rcache_line[5][215].tag_reg.qe       = reg2hw.tag_1495.qe;
  assign rcache_line[5][215].tag_reg.re       = reg2hw.tag_1495.re;
  assign rcache_line[5][215].status_reg.status = reg2hw.status_1495.q;//status_reg_t'(reg2hw.status_1495.q);
  assign rcache_line[5][215].status_reg.qe    = reg2hw.status_1495.qe;
  assign rcache_line[5][215].status_reg.re    = reg2hw.status_1495.re;


  assign rcache_line[5][216].tag_reg.tag      = reg2hw.tag_1496.q;
  assign rcache_line[5][216].tag_reg.qe       = reg2hw.tag_1496.qe;
  assign rcache_line[5][216].tag_reg.re       = reg2hw.tag_1496.re;
  assign rcache_line[5][216].status_reg.status = reg2hw.status_1496.q;//status_reg_t'(reg2hw.status_1496.q);
  assign rcache_line[5][216].status_reg.qe    = reg2hw.status_1496.qe;
  assign rcache_line[5][216].status_reg.re    = reg2hw.status_1496.re;


  assign rcache_line[5][217].tag_reg.tag      = reg2hw.tag_1497.q;
  assign rcache_line[5][217].tag_reg.qe       = reg2hw.tag_1497.qe;
  assign rcache_line[5][217].tag_reg.re       = reg2hw.tag_1497.re;
  assign rcache_line[5][217].status_reg.status = reg2hw.status_1497.q;//status_reg_t'(reg2hw.status_1497.q);
  assign rcache_line[5][217].status_reg.qe    = reg2hw.status_1497.qe;
  assign rcache_line[5][217].status_reg.re    = reg2hw.status_1497.re;


  assign rcache_line[5][218].tag_reg.tag      = reg2hw.tag_1498.q;
  assign rcache_line[5][218].tag_reg.qe       = reg2hw.tag_1498.qe;
  assign rcache_line[5][218].tag_reg.re       = reg2hw.tag_1498.re;
  assign rcache_line[5][218].status_reg.status = reg2hw.status_1498.q;//status_reg_t'(reg2hw.status_1498.q);
  assign rcache_line[5][218].status_reg.qe    = reg2hw.status_1498.qe;
  assign rcache_line[5][218].status_reg.re    = reg2hw.status_1498.re;


  assign rcache_line[5][219].tag_reg.tag      = reg2hw.tag_1499.q;
  assign rcache_line[5][219].tag_reg.qe       = reg2hw.tag_1499.qe;
  assign rcache_line[5][219].tag_reg.re       = reg2hw.tag_1499.re;
  assign rcache_line[5][219].status_reg.status = reg2hw.status_1499.q;//status_reg_t'(reg2hw.status_1499.q);
  assign rcache_line[5][219].status_reg.qe    = reg2hw.status_1499.qe;
  assign rcache_line[5][219].status_reg.re    = reg2hw.status_1499.re;


  assign rcache_line[5][220].tag_reg.tag      = reg2hw.tag_1500.q;
  assign rcache_line[5][220].tag_reg.qe       = reg2hw.tag_1500.qe;
  assign rcache_line[5][220].tag_reg.re       = reg2hw.tag_1500.re;
  assign rcache_line[5][220].status_reg.status = reg2hw.status_1500.q;//status_reg_t'(reg2hw.status_1500.q);
  assign rcache_line[5][220].status_reg.qe    = reg2hw.status_1500.qe;
  assign rcache_line[5][220].status_reg.re    = reg2hw.status_1500.re;


  assign rcache_line[5][221].tag_reg.tag      = reg2hw.tag_1501.q;
  assign rcache_line[5][221].tag_reg.qe       = reg2hw.tag_1501.qe;
  assign rcache_line[5][221].tag_reg.re       = reg2hw.tag_1501.re;
  assign rcache_line[5][221].status_reg.status = reg2hw.status_1501.q;//status_reg_t'(reg2hw.status_1501.q);
  assign rcache_line[5][221].status_reg.qe    = reg2hw.status_1501.qe;
  assign rcache_line[5][221].status_reg.re    = reg2hw.status_1501.re;


  assign rcache_line[5][222].tag_reg.tag      = reg2hw.tag_1502.q;
  assign rcache_line[5][222].tag_reg.qe       = reg2hw.tag_1502.qe;
  assign rcache_line[5][222].tag_reg.re       = reg2hw.tag_1502.re;
  assign rcache_line[5][222].status_reg.status = reg2hw.status_1502.q;//status_reg_t'(reg2hw.status_1502.q);
  assign rcache_line[5][222].status_reg.qe    = reg2hw.status_1502.qe;
  assign rcache_line[5][222].status_reg.re    = reg2hw.status_1502.re;


  assign rcache_line[5][223].tag_reg.tag      = reg2hw.tag_1503.q;
  assign rcache_line[5][223].tag_reg.qe       = reg2hw.tag_1503.qe;
  assign rcache_line[5][223].tag_reg.re       = reg2hw.tag_1503.re;
  assign rcache_line[5][223].status_reg.status = reg2hw.status_1503.q;//status_reg_t'(reg2hw.status_1503.q);
  assign rcache_line[5][223].status_reg.qe    = reg2hw.status_1503.qe;
  assign rcache_line[5][223].status_reg.re    = reg2hw.status_1503.re;


  assign rcache_line[5][224].tag_reg.tag      = reg2hw.tag_1504.q;
  assign rcache_line[5][224].tag_reg.qe       = reg2hw.tag_1504.qe;
  assign rcache_line[5][224].tag_reg.re       = reg2hw.tag_1504.re;
  assign rcache_line[5][224].status_reg.status = reg2hw.status_1504.q;//status_reg_t'(reg2hw.status_1504.q);
  assign rcache_line[5][224].status_reg.qe    = reg2hw.status_1504.qe;
  assign rcache_line[5][224].status_reg.re    = reg2hw.status_1504.re;


  assign rcache_line[5][225].tag_reg.tag      = reg2hw.tag_1505.q;
  assign rcache_line[5][225].tag_reg.qe       = reg2hw.tag_1505.qe;
  assign rcache_line[5][225].tag_reg.re       = reg2hw.tag_1505.re;
  assign rcache_line[5][225].status_reg.status = reg2hw.status_1505.q;//status_reg_t'(reg2hw.status_1505.q);
  assign rcache_line[5][225].status_reg.qe    = reg2hw.status_1505.qe;
  assign rcache_line[5][225].status_reg.re    = reg2hw.status_1505.re;


  assign rcache_line[5][226].tag_reg.tag      = reg2hw.tag_1506.q;
  assign rcache_line[5][226].tag_reg.qe       = reg2hw.tag_1506.qe;
  assign rcache_line[5][226].tag_reg.re       = reg2hw.tag_1506.re;
  assign rcache_line[5][226].status_reg.status = reg2hw.status_1506.q;//status_reg_t'(reg2hw.status_1506.q);
  assign rcache_line[5][226].status_reg.qe    = reg2hw.status_1506.qe;
  assign rcache_line[5][226].status_reg.re    = reg2hw.status_1506.re;


  assign rcache_line[5][227].tag_reg.tag      = reg2hw.tag_1507.q;
  assign rcache_line[5][227].tag_reg.qe       = reg2hw.tag_1507.qe;
  assign rcache_line[5][227].tag_reg.re       = reg2hw.tag_1507.re;
  assign rcache_line[5][227].status_reg.status = reg2hw.status_1507.q;//status_reg_t'(reg2hw.status_1507.q);
  assign rcache_line[5][227].status_reg.qe    = reg2hw.status_1507.qe;
  assign rcache_line[5][227].status_reg.re    = reg2hw.status_1507.re;


  assign rcache_line[5][228].tag_reg.tag      = reg2hw.tag_1508.q;
  assign rcache_line[5][228].tag_reg.qe       = reg2hw.tag_1508.qe;
  assign rcache_line[5][228].tag_reg.re       = reg2hw.tag_1508.re;
  assign rcache_line[5][228].status_reg.status = reg2hw.status_1508.q;//status_reg_t'(reg2hw.status_1508.q);
  assign rcache_line[5][228].status_reg.qe    = reg2hw.status_1508.qe;
  assign rcache_line[5][228].status_reg.re    = reg2hw.status_1508.re;


  assign rcache_line[5][229].tag_reg.tag      = reg2hw.tag_1509.q;
  assign rcache_line[5][229].tag_reg.qe       = reg2hw.tag_1509.qe;
  assign rcache_line[5][229].tag_reg.re       = reg2hw.tag_1509.re;
  assign rcache_line[5][229].status_reg.status = reg2hw.status_1509.q;//status_reg_t'(reg2hw.status_1509.q);
  assign rcache_line[5][229].status_reg.qe    = reg2hw.status_1509.qe;
  assign rcache_line[5][229].status_reg.re    = reg2hw.status_1509.re;


  assign rcache_line[5][230].tag_reg.tag      = reg2hw.tag_1510.q;
  assign rcache_line[5][230].tag_reg.qe       = reg2hw.tag_1510.qe;
  assign rcache_line[5][230].tag_reg.re       = reg2hw.tag_1510.re;
  assign rcache_line[5][230].status_reg.status = reg2hw.status_1510.q;//status_reg_t'(reg2hw.status_1510.q);
  assign rcache_line[5][230].status_reg.qe    = reg2hw.status_1510.qe;
  assign rcache_line[5][230].status_reg.re    = reg2hw.status_1510.re;


  assign rcache_line[5][231].tag_reg.tag      = reg2hw.tag_1511.q;
  assign rcache_line[5][231].tag_reg.qe       = reg2hw.tag_1511.qe;
  assign rcache_line[5][231].tag_reg.re       = reg2hw.tag_1511.re;
  assign rcache_line[5][231].status_reg.status = reg2hw.status_1511.q;//status_reg_t'(reg2hw.status_1511.q);
  assign rcache_line[5][231].status_reg.qe    = reg2hw.status_1511.qe;
  assign rcache_line[5][231].status_reg.re    = reg2hw.status_1511.re;


  assign rcache_line[5][232].tag_reg.tag      = reg2hw.tag_1512.q;
  assign rcache_line[5][232].tag_reg.qe       = reg2hw.tag_1512.qe;
  assign rcache_line[5][232].tag_reg.re       = reg2hw.tag_1512.re;
  assign rcache_line[5][232].status_reg.status = reg2hw.status_1512.q;//status_reg_t'(reg2hw.status_1512.q);
  assign rcache_line[5][232].status_reg.qe    = reg2hw.status_1512.qe;
  assign rcache_line[5][232].status_reg.re    = reg2hw.status_1512.re;


  assign rcache_line[5][233].tag_reg.tag      = reg2hw.tag_1513.q;
  assign rcache_line[5][233].tag_reg.qe       = reg2hw.tag_1513.qe;
  assign rcache_line[5][233].tag_reg.re       = reg2hw.tag_1513.re;
  assign rcache_line[5][233].status_reg.status = reg2hw.status_1513.q;//status_reg_t'(reg2hw.status_1513.q);
  assign rcache_line[5][233].status_reg.qe    = reg2hw.status_1513.qe;
  assign rcache_line[5][233].status_reg.re    = reg2hw.status_1513.re;


  assign rcache_line[5][234].tag_reg.tag      = reg2hw.tag_1514.q;
  assign rcache_line[5][234].tag_reg.qe       = reg2hw.tag_1514.qe;
  assign rcache_line[5][234].tag_reg.re       = reg2hw.tag_1514.re;
  assign rcache_line[5][234].status_reg.status = reg2hw.status_1514.q;//status_reg_t'(reg2hw.status_1514.q);
  assign rcache_line[5][234].status_reg.qe    = reg2hw.status_1514.qe;
  assign rcache_line[5][234].status_reg.re    = reg2hw.status_1514.re;


  assign rcache_line[5][235].tag_reg.tag      = reg2hw.tag_1515.q;
  assign rcache_line[5][235].tag_reg.qe       = reg2hw.tag_1515.qe;
  assign rcache_line[5][235].tag_reg.re       = reg2hw.tag_1515.re;
  assign rcache_line[5][235].status_reg.status = reg2hw.status_1515.q;//status_reg_t'(reg2hw.status_1515.q);
  assign rcache_line[5][235].status_reg.qe    = reg2hw.status_1515.qe;
  assign rcache_line[5][235].status_reg.re    = reg2hw.status_1515.re;


  assign rcache_line[5][236].tag_reg.tag      = reg2hw.tag_1516.q;
  assign rcache_line[5][236].tag_reg.qe       = reg2hw.tag_1516.qe;
  assign rcache_line[5][236].tag_reg.re       = reg2hw.tag_1516.re;
  assign rcache_line[5][236].status_reg.status = reg2hw.status_1516.q;//status_reg_t'(reg2hw.status_1516.q);
  assign rcache_line[5][236].status_reg.qe    = reg2hw.status_1516.qe;
  assign rcache_line[5][236].status_reg.re    = reg2hw.status_1516.re;


  assign rcache_line[5][237].tag_reg.tag      = reg2hw.tag_1517.q;
  assign rcache_line[5][237].tag_reg.qe       = reg2hw.tag_1517.qe;
  assign rcache_line[5][237].tag_reg.re       = reg2hw.tag_1517.re;
  assign rcache_line[5][237].status_reg.status = reg2hw.status_1517.q;//status_reg_t'(reg2hw.status_1517.q);
  assign rcache_line[5][237].status_reg.qe    = reg2hw.status_1517.qe;
  assign rcache_line[5][237].status_reg.re    = reg2hw.status_1517.re;


  assign rcache_line[5][238].tag_reg.tag      = reg2hw.tag_1518.q;
  assign rcache_line[5][238].tag_reg.qe       = reg2hw.tag_1518.qe;
  assign rcache_line[5][238].tag_reg.re       = reg2hw.tag_1518.re;
  assign rcache_line[5][238].status_reg.status = reg2hw.status_1518.q;//status_reg_t'(reg2hw.status_1518.q);
  assign rcache_line[5][238].status_reg.qe    = reg2hw.status_1518.qe;
  assign rcache_line[5][238].status_reg.re    = reg2hw.status_1518.re;


  assign rcache_line[5][239].tag_reg.tag      = reg2hw.tag_1519.q;
  assign rcache_line[5][239].tag_reg.qe       = reg2hw.tag_1519.qe;
  assign rcache_line[5][239].tag_reg.re       = reg2hw.tag_1519.re;
  assign rcache_line[5][239].status_reg.status = reg2hw.status_1519.q;//status_reg_t'(reg2hw.status_1519.q);
  assign rcache_line[5][239].status_reg.qe    = reg2hw.status_1519.qe;
  assign rcache_line[5][239].status_reg.re    = reg2hw.status_1519.re;


  assign rcache_line[5][240].tag_reg.tag      = reg2hw.tag_1520.q;
  assign rcache_line[5][240].tag_reg.qe       = reg2hw.tag_1520.qe;
  assign rcache_line[5][240].tag_reg.re       = reg2hw.tag_1520.re;
  assign rcache_line[5][240].status_reg.status = reg2hw.status_1520.q;//status_reg_t'(reg2hw.status_1520.q);
  assign rcache_line[5][240].status_reg.qe    = reg2hw.status_1520.qe;
  assign rcache_line[5][240].status_reg.re    = reg2hw.status_1520.re;


  assign rcache_line[5][241].tag_reg.tag      = reg2hw.tag_1521.q;
  assign rcache_line[5][241].tag_reg.qe       = reg2hw.tag_1521.qe;
  assign rcache_line[5][241].tag_reg.re       = reg2hw.tag_1521.re;
  assign rcache_line[5][241].status_reg.status = reg2hw.status_1521.q;//status_reg_t'(reg2hw.status_1521.q);
  assign rcache_line[5][241].status_reg.qe    = reg2hw.status_1521.qe;
  assign rcache_line[5][241].status_reg.re    = reg2hw.status_1521.re;


  assign rcache_line[5][242].tag_reg.tag      = reg2hw.tag_1522.q;
  assign rcache_line[5][242].tag_reg.qe       = reg2hw.tag_1522.qe;
  assign rcache_line[5][242].tag_reg.re       = reg2hw.tag_1522.re;
  assign rcache_line[5][242].status_reg.status = reg2hw.status_1522.q;//status_reg_t'(reg2hw.status_1522.q);
  assign rcache_line[5][242].status_reg.qe    = reg2hw.status_1522.qe;
  assign rcache_line[5][242].status_reg.re    = reg2hw.status_1522.re;


  assign rcache_line[5][243].tag_reg.tag      = reg2hw.tag_1523.q;
  assign rcache_line[5][243].tag_reg.qe       = reg2hw.tag_1523.qe;
  assign rcache_line[5][243].tag_reg.re       = reg2hw.tag_1523.re;
  assign rcache_line[5][243].status_reg.status = reg2hw.status_1523.q;//status_reg_t'(reg2hw.status_1523.q);
  assign rcache_line[5][243].status_reg.qe    = reg2hw.status_1523.qe;
  assign rcache_line[5][243].status_reg.re    = reg2hw.status_1523.re;


  assign rcache_line[5][244].tag_reg.tag      = reg2hw.tag_1524.q;
  assign rcache_line[5][244].tag_reg.qe       = reg2hw.tag_1524.qe;
  assign rcache_line[5][244].tag_reg.re       = reg2hw.tag_1524.re;
  assign rcache_line[5][244].status_reg.status = reg2hw.status_1524.q;//status_reg_t'(reg2hw.status_1524.q);
  assign rcache_line[5][244].status_reg.qe    = reg2hw.status_1524.qe;
  assign rcache_line[5][244].status_reg.re    = reg2hw.status_1524.re;


  assign rcache_line[5][245].tag_reg.tag      = reg2hw.tag_1525.q;
  assign rcache_line[5][245].tag_reg.qe       = reg2hw.tag_1525.qe;
  assign rcache_line[5][245].tag_reg.re       = reg2hw.tag_1525.re;
  assign rcache_line[5][245].status_reg.status = reg2hw.status_1525.q;//status_reg_t'(reg2hw.status_1525.q);
  assign rcache_line[5][245].status_reg.qe    = reg2hw.status_1525.qe;
  assign rcache_line[5][245].status_reg.re    = reg2hw.status_1525.re;


  assign rcache_line[5][246].tag_reg.tag      = reg2hw.tag_1526.q;
  assign rcache_line[5][246].tag_reg.qe       = reg2hw.tag_1526.qe;
  assign rcache_line[5][246].tag_reg.re       = reg2hw.tag_1526.re;
  assign rcache_line[5][246].status_reg.status = reg2hw.status_1526.q;//status_reg_t'(reg2hw.status_1526.q);
  assign rcache_line[5][246].status_reg.qe    = reg2hw.status_1526.qe;
  assign rcache_line[5][246].status_reg.re    = reg2hw.status_1526.re;


  assign rcache_line[5][247].tag_reg.tag      = reg2hw.tag_1527.q;
  assign rcache_line[5][247].tag_reg.qe       = reg2hw.tag_1527.qe;
  assign rcache_line[5][247].tag_reg.re       = reg2hw.tag_1527.re;
  assign rcache_line[5][247].status_reg.status = reg2hw.status_1527.q;//status_reg_t'(reg2hw.status_1527.q);
  assign rcache_line[5][247].status_reg.qe    = reg2hw.status_1527.qe;
  assign rcache_line[5][247].status_reg.re    = reg2hw.status_1527.re;


  assign rcache_line[5][248].tag_reg.tag      = reg2hw.tag_1528.q;
  assign rcache_line[5][248].tag_reg.qe       = reg2hw.tag_1528.qe;
  assign rcache_line[5][248].tag_reg.re       = reg2hw.tag_1528.re;
  assign rcache_line[5][248].status_reg.status = reg2hw.status_1528.q;//status_reg_t'(reg2hw.status_1528.q);
  assign rcache_line[5][248].status_reg.qe    = reg2hw.status_1528.qe;
  assign rcache_line[5][248].status_reg.re    = reg2hw.status_1528.re;


  assign rcache_line[5][249].tag_reg.tag      = reg2hw.tag_1529.q;
  assign rcache_line[5][249].tag_reg.qe       = reg2hw.tag_1529.qe;
  assign rcache_line[5][249].tag_reg.re       = reg2hw.tag_1529.re;
  assign rcache_line[5][249].status_reg.status = reg2hw.status_1529.q;//status_reg_t'(reg2hw.status_1529.q);
  assign rcache_line[5][249].status_reg.qe    = reg2hw.status_1529.qe;
  assign rcache_line[5][249].status_reg.re    = reg2hw.status_1529.re;


  assign rcache_line[5][250].tag_reg.tag      = reg2hw.tag_1530.q;
  assign rcache_line[5][250].tag_reg.qe       = reg2hw.tag_1530.qe;
  assign rcache_line[5][250].tag_reg.re       = reg2hw.tag_1530.re;
  assign rcache_line[5][250].status_reg.status = reg2hw.status_1530.q;//status_reg_t'(reg2hw.status_1530.q);
  assign rcache_line[5][250].status_reg.qe    = reg2hw.status_1530.qe;
  assign rcache_line[5][250].status_reg.re    = reg2hw.status_1530.re;


  assign rcache_line[5][251].tag_reg.tag      = reg2hw.tag_1531.q;
  assign rcache_line[5][251].tag_reg.qe       = reg2hw.tag_1531.qe;
  assign rcache_line[5][251].tag_reg.re       = reg2hw.tag_1531.re;
  assign rcache_line[5][251].status_reg.status = reg2hw.status_1531.q;//status_reg_t'(reg2hw.status_1531.q);
  assign rcache_line[5][251].status_reg.qe    = reg2hw.status_1531.qe;
  assign rcache_line[5][251].status_reg.re    = reg2hw.status_1531.re;


  assign rcache_line[5][252].tag_reg.tag      = reg2hw.tag_1532.q;
  assign rcache_line[5][252].tag_reg.qe       = reg2hw.tag_1532.qe;
  assign rcache_line[5][252].tag_reg.re       = reg2hw.tag_1532.re;
  assign rcache_line[5][252].status_reg.status = reg2hw.status_1532.q;//status_reg_t'(reg2hw.status_1532.q);
  assign rcache_line[5][252].status_reg.qe    = reg2hw.status_1532.qe;
  assign rcache_line[5][252].status_reg.re    = reg2hw.status_1532.re;


  assign rcache_line[5][253].tag_reg.tag      = reg2hw.tag_1533.q;
  assign rcache_line[5][253].tag_reg.qe       = reg2hw.tag_1533.qe;
  assign rcache_line[5][253].tag_reg.re       = reg2hw.tag_1533.re;
  assign rcache_line[5][253].status_reg.status = reg2hw.status_1533.q;//status_reg_t'(reg2hw.status_1533.q);
  assign rcache_line[5][253].status_reg.qe    = reg2hw.status_1533.qe;
  assign rcache_line[5][253].status_reg.re    = reg2hw.status_1533.re;


  assign rcache_line[5][254].tag_reg.tag      = reg2hw.tag_1534.q;
  assign rcache_line[5][254].tag_reg.qe       = reg2hw.tag_1534.qe;
  assign rcache_line[5][254].tag_reg.re       = reg2hw.tag_1534.re;
  assign rcache_line[5][254].status_reg.status = reg2hw.status_1534.q;//status_reg_t'(reg2hw.status_1534.q);
  assign rcache_line[5][254].status_reg.qe    = reg2hw.status_1534.qe;
  assign rcache_line[5][254].status_reg.re    = reg2hw.status_1534.re;


  assign rcache_line[5][255].tag_reg.tag      = reg2hw.tag_1535.q;
  assign rcache_line[5][255].tag_reg.qe       = reg2hw.tag_1535.qe;
  assign rcache_line[5][255].tag_reg.re       = reg2hw.tag_1535.re;
  assign rcache_line[5][255].status_reg.status = reg2hw.status_1535.q;//status_reg_t'(reg2hw.status_1535.q);
  assign rcache_line[5][255].status_reg.qe    = reg2hw.status_1535.qe;
  assign rcache_line[5][255].status_reg.re    = reg2hw.status_1535.re;


  assign rcache_line[6][0].tag_reg.tag      = reg2hw.tag_1536.q;
  assign rcache_line[6][0].tag_reg.qe       = reg2hw.tag_1536.qe;
  assign rcache_line[6][0].tag_reg.re       = reg2hw.tag_1536.re;
  assign rcache_line[6][0].status_reg.status = reg2hw.status_1536.q;//status_reg_t'(reg2hw.status_1536.q);
  assign rcache_line[6][0].status_reg.qe    = reg2hw.status_1536.qe;
  assign rcache_line[6][0].status_reg.re    = reg2hw.status_1536.re;


  assign rcache_line[6][1].tag_reg.tag      = reg2hw.tag_1537.q;
  assign rcache_line[6][1].tag_reg.qe       = reg2hw.tag_1537.qe;
  assign rcache_line[6][1].tag_reg.re       = reg2hw.tag_1537.re;
  assign rcache_line[6][1].status_reg.status = reg2hw.status_1537.q;//status_reg_t'(reg2hw.status_1537.q);
  assign rcache_line[6][1].status_reg.qe    = reg2hw.status_1537.qe;
  assign rcache_line[6][1].status_reg.re    = reg2hw.status_1537.re;


  assign rcache_line[6][2].tag_reg.tag      = reg2hw.tag_1538.q;
  assign rcache_line[6][2].tag_reg.qe       = reg2hw.tag_1538.qe;
  assign rcache_line[6][2].tag_reg.re       = reg2hw.tag_1538.re;
  assign rcache_line[6][2].status_reg.status = reg2hw.status_1538.q;//status_reg_t'(reg2hw.status_1538.q);
  assign rcache_line[6][2].status_reg.qe    = reg2hw.status_1538.qe;
  assign rcache_line[6][2].status_reg.re    = reg2hw.status_1538.re;


  assign rcache_line[6][3].tag_reg.tag      = reg2hw.tag_1539.q;
  assign rcache_line[6][3].tag_reg.qe       = reg2hw.tag_1539.qe;
  assign rcache_line[6][3].tag_reg.re       = reg2hw.tag_1539.re;
  assign rcache_line[6][3].status_reg.status = reg2hw.status_1539.q;//status_reg_t'(reg2hw.status_1539.q);
  assign rcache_line[6][3].status_reg.qe    = reg2hw.status_1539.qe;
  assign rcache_line[6][3].status_reg.re    = reg2hw.status_1539.re;


  assign rcache_line[6][4].tag_reg.tag      = reg2hw.tag_1540.q;
  assign rcache_line[6][4].tag_reg.qe       = reg2hw.tag_1540.qe;
  assign rcache_line[6][4].tag_reg.re       = reg2hw.tag_1540.re;
  assign rcache_line[6][4].status_reg.status = reg2hw.status_1540.q;//status_reg_t'(reg2hw.status_1540.q);
  assign rcache_line[6][4].status_reg.qe    = reg2hw.status_1540.qe;
  assign rcache_line[6][4].status_reg.re    = reg2hw.status_1540.re;


  assign rcache_line[6][5].tag_reg.tag      = reg2hw.tag_1541.q;
  assign rcache_line[6][5].tag_reg.qe       = reg2hw.tag_1541.qe;
  assign rcache_line[6][5].tag_reg.re       = reg2hw.tag_1541.re;
  assign rcache_line[6][5].status_reg.status = reg2hw.status_1541.q;//status_reg_t'(reg2hw.status_1541.q);
  assign rcache_line[6][5].status_reg.qe    = reg2hw.status_1541.qe;
  assign rcache_line[6][5].status_reg.re    = reg2hw.status_1541.re;


  assign rcache_line[6][6].tag_reg.tag      = reg2hw.tag_1542.q;
  assign rcache_line[6][6].tag_reg.qe       = reg2hw.tag_1542.qe;
  assign rcache_line[6][6].tag_reg.re       = reg2hw.tag_1542.re;
  assign rcache_line[6][6].status_reg.status = reg2hw.status_1542.q;//status_reg_t'(reg2hw.status_1542.q);
  assign rcache_line[6][6].status_reg.qe    = reg2hw.status_1542.qe;
  assign rcache_line[6][6].status_reg.re    = reg2hw.status_1542.re;


  assign rcache_line[6][7].tag_reg.tag      = reg2hw.tag_1543.q;
  assign rcache_line[6][7].tag_reg.qe       = reg2hw.tag_1543.qe;
  assign rcache_line[6][7].tag_reg.re       = reg2hw.tag_1543.re;
  assign rcache_line[6][7].status_reg.status = reg2hw.status_1543.q;//status_reg_t'(reg2hw.status_1543.q);
  assign rcache_line[6][7].status_reg.qe    = reg2hw.status_1543.qe;
  assign rcache_line[6][7].status_reg.re    = reg2hw.status_1543.re;


  assign rcache_line[6][8].tag_reg.tag      = reg2hw.tag_1544.q;
  assign rcache_line[6][8].tag_reg.qe       = reg2hw.tag_1544.qe;
  assign rcache_line[6][8].tag_reg.re       = reg2hw.tag_1544.re;
  assign rcache_line[6][8].status_reg.status = reg2hw.status_1544.q;//status_reg_t'(reg2hw.status_1544.q);
  assign rcache_line[6][8].status_reg.qe    = reg2hw.status_1544.qe;
  assign rcache_line[6][8].status_reg.re    = reg2hw.status_1544.re;


  assign rcache_line[6][9].tag_reg.tag      = reg2hw.tag_1545.q;
  assign rcache_line[6][9].tag_reg.qe       = reg2hw.tag_1545.qe;
  assign rcache_line[6][9].tag_reg.re       = reg2hw.tag_1545.re;
  assign rcache_line[6][9].status_reg.status = reg2hw.status_1545.q;//status_reg_t'(reg2hw.status_1545.q);
  assign rcache_line[6][9].status_reg.qe    = reg2hw.status_1545.qe;
  assign rcache_line[6][9].status_reg.re    = reg2hw.status_1545.re;


  assign rcache_line[6][10].tag_reg.tag      = reg2hw.tag_1546.q;
  assign rcache_line[6][10].tag_reg.qe       = reg2hw.tag_1546.qe;
  assign rcache_line[6][10].tag_reg.re       = reg2hw.tag_1546.re;
  assign rcache_line[6][10].status_reg.status = reg2hw.status_1546.q;//status_reg_t'(reg2hw.status_1546.q);
  assign rcache_line[6][10].status_reg.qe    = reg2hw.status_1546.qe;
  assign rcache_line[6][10].status_reg.re    = reg2hw.status_1546.re;


  assign rcache_line[6][11].tag_reg.tag      = reg2hw.tag_1547.q;
  assign rcache_line[6][11].tag_reg.qe       = reg2hw.tag_1547.qe;
  assign rcache_line[6][11].tag_reg.re       = reg2hw.tag_1547.re;
  assign rcache_line[6][11].status_reg.status = reg2hw.status_1547.q;//status_reg_t'(reg2hw.status_1547.q);
  assign rcache_line[6][11].status_reg.qe    = reg2hw.status_1547.qe;
  assign rcache_line[6][11].status_reg.re    = reg2hw.status_1547.re;


  assign rcache_line[6][12].tag_reg.tag      = reg2hw.tag_1548.q;
  assign rcache_line[6][12].tag_reg.qe       = reg2hw.tag_1548.qe;
  assign rcache_line[6][12].tag_reg.re       = reg2hw.tag_1548.re;
  assign rcache_line[6][12].status_reg.status = reg2hw.status_1548.q;//status_reg_t'(reg2hw.status_1548.q);
  assign rcache_line[6][12].status_reg.qe    = reg2hw.status_1548.qe;
  assign rcache_line[6][12].status_reg.re    = reg2hw.status_1548.re;


  assign rcache_line[6][13].tag_reg.tag      = reg2hw.tag_1549.q;
  assign rcache_line[6][13].tag_reg.qe       = reg2hw.tag_1549.qe;
  assign rcache_line[6][13].tag_reg.re       = reg2hw.tag_1549.re;
  assign rcache_line[6][13].status_reg.status = reg2hw.status_1549.q;//status_reg_t'(reg2hw.status_1549.q);
  assign rcache_line[6][13].status_reg.qe    = reg2hw.status_1549.qe;
  assign rcache_line[6][13].status_reg.re    = reg2hw.status_1549.re;


  assign rcache_line[6][14].tag_reg.tag      = reg2hw.tag_1550.q;
  assign rcache_line[6][14].tag_reg.qe       = reg2hw.tag_1550.qe;
  assign rcache_line[6][14].tag_reg.re       = reg2hw.tag_1550.re;
  assign rcache_line[6][14].status_reg.status = reg2hw.status_1550.q;//status_reg_t'(reg2hw.status_1550.q);
  assign rcache_line[6][14].status_reg.qe    = reg2hw.status_1550.qe;
  assign rcache_line[6][14].status_reg.re    = reg2hw.status_1550.re;


  assign rcache_line[6][15].tag_reg.tag      = reg2hw.tag_1551.q;
  assign rcache_line[6][15].tag_reg.qe       = reg2hw.tag_1551.qe;
  assign rcache_line[6][15].tag_reg.re       = reg2hw.tag_1551.re;
  assign rcache_line[6][15].status_reg.status = reg2hw.status_1551.q;//status_reg_t'(reg2hw.status_1551.q);
  assign rcache_line[6][15].status_reg.qe    = reg2hw.status_1551.qe;
  assign rcache_line[6][15].status_reg.re    = reg2hw.status_1551.re;


  assign rcache_line[6][16].tag_reg.tag      = reg2hw.tag_1552.q;
  assign rcache_line[6][16].tag_reg.qe       = reg2hw.tag_1552.qe;
  assign rcache_line[6][16].tag_reg.re       = reg2hw.tag_1552.re;
  assign rcache_line[6][16].status_reg.status = reg2hw.status_1552.q;//status_reg_t'(reg2hw.status_1552.q);
  assign rcache_line[6][16].status_reg.qe    = reg2hw.status_1552.qe;
  assign rcache_line[6][16].status_reg.re    = reg2hw.status_1552.re;


  assign rcache_line[6][17].tag_reg.tag      = reg2hw.tag_1553.q;
  assign rcache_line[6][17].tag_reg.qe       = reg2hw.tag_1553.qe;
  assign rcache_line[6][17].tag_reg.re       = reg2hw.tag_1553.re;
  assign rcache_line[6][17].status_reg.status = reg2hw.status_1553.q;//status_reg_t'(reg2hw.status_1553.q);
  assign rcache_line[6][17].status_reg.qe    = reg2hw.status_1553.qe;
  assign rcache_line[6][17].status_reg.re    = reg2hw.status_1553.re;


  assign rcache_line[6][18].tag_reg.tag      = reg2hw.tag_1554.q;
  assign rcache_line[6][18].tag_reg.qe       = reg2hw.tag_1554.qe;
  assign rcache_line[6][18].tag_reg.re       = reg2hw.tag_1554.re;
  assign rcache_line[6][18].status_reg.status = reg2hw.status_1554.q;//status_reg_t'(reg2hw.status_1554.q);
  assign rcache_line[6][18].status_reg.qe    = reg2hw.status_1554.qe;
  assign rcache_line[6][18].status_reg.re    = reg2hw.status_1554.re;


  assign rcache_line[6][19].tag_reg.tag      = reg2hw.tag_1555.q;
  assign rcache_line[6][19].tag_reg.qe       = reg2hw.tag_1555.qe;
  assign rcache_line[6][19].tag_reg.re       = reg2hw.tag_1555.re;
  assign rcache_line[6][19].status_reg.status = reg2hw.status_1555.q;//status_reg_t'(reg2hw.status_1555.q);
  assign rcache_line[6][19].status_reg.qe    = reg2hw.status_1555.qe;
  assign rcache_line[6][19].status_reg.re    = reg2hw.status_1555.re;


  assign rcache_line[6][20].tag_reg.tag      = reg2hw.tag_1556.q;
  assign rcache_line[6][20].tag_reg.qe       = reg2hw.tag_1556.qe;
  assign rcache_line[6][20].tag_reg.re       = reg2hw.tag_1556.re;
  assign rcache_line[6][20].status_reg.status = reg2hw.status_1556.q;//status_reg_t'(reg2hw.status_1556.q);
  assign rcache_line[6][20].status_reg.qe    = reg2hw.status_1556.qe;
  assign rcache_line[6][20].status_reg.re    = reg2hw.status_1556.re;


  assign rcache_line[6][21].tag_reg.tag      = reg2hw.tag_1557.q;
  assign rcache_line[6][21].tag_reg.qe       = reg2hw.tag_1557.qe;
  assign rcache_line[6][21].tag_reg.re       = reg2hw.tag_1557.re;
  assign rcache_line[6][21].status_reg.status = reg2hw.status_1557.q;//status_reg_t'(reg2hw.status_1557.q);
  assign rcache_line[6][21].status_reg.qe    = reg2hw.status_1557.qe;
  assign rcache_line[6][21].status_reg.re    = reg2hw.status_1557.re;


  assign rcache_line[6][22].tag_reg.tag      = reg2hw.tag_1558.q;
  assign rcache_line[6][22].tag_reg.qe       = reg2hw.tag_1558.qe;
  assign rcache_line[6][22].tag_reg.re       = reg2hw.tag_1558.re;
  assign rcache_line[6][22].status_reg.status = reg2hw.status_1558.q;//status_reg_t'(reg2hw.status_1558.q);
  assign rcache_line[6][22].status_reg.qe    = reg2hw.status_1558.qe;
  assign rcache_line[6][22].status_reg.re    = reg2hw.status_1558.re;


  assign rcache_line[6][23].tag_reg.tag      = reg2hw.tag_1559.q;
  assign rcache_line[6][23].tag_reg.qe       = reg2hw.tag_1559.qe;
  assign rcache_line[6][23].tag_reg.re       = reg2hw.tag_1559.re;
  assign rcache_line[6][23].status_reg.status = reg2hw.status_1559.q;//status_reg_t'(reg2hw.status_1559.q);
  assign rcache_line[6][23].status_reg.qe    = reg2hw.status_1559.qe;
  assign rcache_line[6][23].status_reg.re    = reg2hw.status_1559.re;


  assign rcache_line[6][24].tag_reg.tag      = reg2hw.tag_1560.q;
  assign rcache_line[6][24].tag_reg.qe       = reg2hw.tag_1560.qe;
  assign rcache_line[6][24].tag_reg.re       = reg2hw.tag_1560.re;
  assign rcache_line[6][24].status_reg.status = reg2hw.status_1560.q;//status_reg_t'(reg2hw.status_1560.q);
  assign rcache_line[6][24].status_reg.qe    = reg2hw.status_1560.qe;
  assign rcache_line[6][24].status_reg.re    = reg2hw.status_1560.re;


  assign rcache_line[6][25].tag_reg.tag      = reg2hw.tag_1561.q;
  assign rcache_line[6][25].tag_reg.qe       = reg2hw.tag_1561.qe;
  assign rcache_line[6][25].tag_reg.re       = reg2hw.tag_1561.re;
  assign rcache_line[6][25].status_reg.status = reg2hw.status_1561.q;//status_reg_t'(reg2hw.status_1561.q);
  assign rcache_line[6][25].status_reg.qe    = reg2hw.status_1561.qe;
  assign rcache_line[6][25].status_reg.re    = reg2hw.status_1561.re;


  assign rcache_line[6][26].tag_reg.tag      = reg2hw.tag_1562.q;
  assign rcache_line[6][26].tag_reg.qe       = reg2hw.tag_1562.qe;
  assign rcache_line[6][26].tag_reg.re       = reg2hw.tag_1562.re;
  assign rcache_line[6][26].status_reg.status = reg2hw.status_1562.q;//status_reg_t'(reg2hw.status_1562.q);
  assign rcache_line[6][26].status_reg.qe    = reg2hw.status_1562.qe;
  assign rcache_line[6][26].status_reg.re    = reg2hw.status_1562.re;


  assign rcache_line[6][27].tag_reg.tag      = reg2hw.tag_1563.q;
  assign rcache_line[6][27].tag_reg.qe       = reg2hw.tag_1563.qe;
  assign rcache_line[6][27].tag_reg.re       = reg2hw.tag_1563.re;
  assign rcache_line[6][27].status_reg.status = reg2hw.status_1563.q;//status_reg_t'(reg2hw.status_1563.q);
  assign rcache_line[6][27].status_reg.qe    = reg2hw.status_1563.qe;
  assign rcache_line[6][27].status_reg.re    = reg2hw.status_1563.re;


  assign rcache_line[6][28].tag_reg.tag      = reg2hw.tag_1564.q;
  assign rcache_line[6][28].tag_reg.qe       = reg2hw.tag_1564.qe;
  assign rcache_line[6][28].tag_reg.re       = reg2hw.tag_1564.re;
  assign rcache_line[6][28].status_reg.status = reg2hw.status_1564.q;//status_reg_t'(reg2hw.status_1564.q);
  assign rcache_line[6][28].status_reg.qe    = reg2hw.status_1564.qe;
  assign rcache_line[6][28].status_reg.re    = reg2hw.status_1564.re;


  assign rcache_line[6][29].tag_reg.tag      = reg2hw.tag_1565.q;
  assign rcache_line[6][29].tag_reg.qe       = reg2hw.tag_1565.qe;
  assign rcache_line[6][29].tag_reg.re       = reg2hw.tag_1565.re;
  assign rcache_line[6][29].status_reg.status = reg2hw.status_1565.q;//status_reg_t'(reg2hw.status_1565.q);
  assign rcache_line[6][29].status_reg.qe    = reg2hw.status_1565.qe;
  assign rcache_line[6][29].status_reg.re    = reg2hw.status_1565.re;


  assign rcache_line[6][30].tag_reg.tag      = reg2hw.tag_1566.q;
  assign rcache_line[6][30].tag_reg.qe       = reg2hw.tag_1566.qe;
  assign rcache_line[6][30].tag_reg.re       = reg2hw.tag_1566.re;
  assign rcache_line[6][30].status_reg.status = reg2hw.status_1566.q;//status_reg_t'(reg2hw.status_1566.q);
  assign rcache_line[6][30].status_reg.qe    = reg2hw.status_1566.qe;
  assign rcache_line[6][30].status_reg.re    = reg2hw.status_1566.re;


  assign rcache_line[6][31].tag_reg.tag      = reg2hw.tag_1567.q;
  assign rcache_line[6][31].tag_reg.qe       = reg2hw.tag_1567.qe;
  assign rcache_line[6][31].tag_reg.re       = reg2hw.tag_1567.re;
  assign rcache_line[6][31].status_reg.status = reg2hw.status_1567.q;//status_reg_t'(reg2hw.status_1567.q);
  assign rcache_line[6][31].status_reg.qe    = reg2hw.status_1567.qe;
  assign rcache_line[6][31].status_reg.re    = reg2hw.status_1567.re;


  assign rcache_line[6][32].tag_reg.tag      = reg2hw.tag_1568.q;
  assign rcache_line[6][32].tag_reg.qe       = reg2hw.tag_1568.qe;
  assign rcache_line[6][32].tag_reg.re       = reg2hw.tag_1568.re;
  assign rcache_line[6][32].status_reg.status = reg2hw.status_1568.q;//status_reg_t'(reg2hw.status_1568.q);
  assign rcache_line[6][32].status_reg.qe    = reg2hw.status_1568.qe;
  assign rcache_line[6][32].status_reg.re    = reg2hw.status_1568.re;


  assign rcache_line[6][33].tag_reg.tag      = reg2hw.tag_1569.q;
  assign rcache_line[6][33].tag_reg.qe       = reg2hw.tag_1569.qe;
  assign rcache_line[6][33].tag_reg.re       = reg2hw.tag_1569.re;
  assign rcache_line[6][33].status_reg.status = reg2hw.status_1569.q;//status_reg_t'(reg2hw.status_1569.q);
  assign rcache_line[6][33].status_reg.qe    = reg2hw.status_1569.qe;
  assign rcache_line[6][33].status_reg.re    = reg2hw.status_1569.re;


  assign rcache_line[6][34].tag_reg.tag      = reg2hw.tag_1570.q;
  assign rcache_line[6][34].tag_reg.qe       = reg2hw.tag_1570.qe;
  assign rcache_line[6][34].tag_reg.re       = reg2hw.tag_1570.re;
  assign rcache_line[6][34].status_reg.status = reg2hw.status_1570.q;//status_reg_t'(reg2hw.status_1570.q);
  assign rcache_line[6][34].status_reg.qe    = reg2hw.status_1570.qe;
  assign rcache_line[6][34].status_reg.re    = reg2hw.status_1570.re;


  assign rcache_line[6][35].tag_reg.tag      = reg2hw.tag_1571.q;
  assign rcache_line[6][35].tag_reg.qe       = reg2hw.tag_1571.qe;
  assign rcache_line[6][35].tag_reg.re       = reg2hw.tag_1571.re;
  assign rcache_line[6][35].status_reg.status = reg2hw.status_1571.q;//status_reg_t'(reg2hw.status_1571.q);
  assign rcache_line[6][35].status_reg.qe    = reg2hw.status_1571.qe;
  assign rcache_line[6][35].status_reg.re    = reg2hw.status_1571.re;


  assign rcache_line[6][36].tag_reg.tag      = reg2hw.tag_1572.q;
  assign rcache_line[6][36].tag_reg.qe       = reg2hw.tag_1572.qe;
  assign rcache_line[6][36].tag_reg.re       = reg2hw.tag_1572.re;
  assign rcache_line[6][36].status_reg.status = reg2hw.status_1572.q;//status_reg_t'(reg2hw.status_1572.q);
  assign rcache_line[6][36].status_reg.qe    = reg2hw.status_1572.qe;
  assign rcache_line[6][36].status_reg.re    = reg2hw.status_1572.re;


  assign rcache_line[6][37].tag_reg.tag      = reg2hw.tag_1573.q;
  assign rcache_line[6][37].tag_reg.qe       = reg2hw.tag_1573.qe;
  assign rcache_line[6][37].tag_reg.re       = reg2hw.tag_1573.re;
  assign rcache_line[6][37].status_reg.status = reg2hw.status_1573.q;//status_reg_t'(reg2hw.status_1573.q);
  assign rcache_line[6][37].status_reg.qe    = reg2hw.status_1573.qe;
  assign rcache_line[6][37].status_reg.re    = reg2hw.status_1573.re;


  assign rcache_line[6][38].tag_reg.tag      = reg2hw.tag_1574.q;
  assign rcache_line[6][38].tag_reg.qe       = reg2hw.tag_1574.qe;
  assign rcache_line[6][38].tag_reg.re       = reg2hw.tag_1574.re;
  assign rcache_line[6][38].status_reg.status = reg2hw.status_1574.q;//status_reg_t'(reg2hw.status_1574.q);
  assign rcache_line[6][38].status_reg.qe    = reg2hw.status_1574.qe;
  assign rcache_line[6][38].status_reg.re    = reg2hw.status_1574.re;


  assign rcache_line[6][39].tag_reg.tag      = reg2hw.tag_1575.q;
  assign rcache_line[6][39].tag_reg.qe       = reg2hw.tag_1575.qe;
  assign rcache_line[6][39].tag_reg.re       = reg2hw.tag_1575.re;
  assign rcache_line[6][39].status_reg.status = reg2hw.status_1575.q;//status_reg_t'(reg2hw.status_1575.q);
  assign rcache_line[6][39].status_reg.qe    = reg2hw.status_1575.qe;
  assign rcache_line[6][39].status_reg.re    = reg2hw.status_1575.re;


  assign rcache_line[6][40].tag_reg.tag      = reg2hw.tag_1576.q;
  assign rcache_line[6][40].tag_reg.qe       = reg2hw.tag_1576.qe;
  assign rcache_line[6][40].tag_reg.re       = reg2hw.tag_1576.re;
  assign rcache_line[6][40].status_reg.status = reg2hw.status_1576.q;//status_reg_t'(reg2hw.status_1576.q);
  assign rcache_line[6][40].status_reg.qe    = reg2hw.status_1576.qe;
  assign rcache_line[6][40].status_reg.re    = reg2hw.status_1576.re;


  assign rcache_line[6][41].tag_reg.tag      = reg2hw.tag_1577.q;
  assign rcache_line[6][41].tag_reg.qe       = reg2hw.tag_1577.qe;
  assign rcache_line[6][41].tag_reg.re       = reg2hw.tag_1577.re;
  assign rcache_line[6][41].status_reg.status = reg2hw.status_1577.q;//status_reg_t'(reg2hw.status_1577.q);
  assign rcache_line[6][41].status_reg.qe    = reg2hw.status_1577.qe;
  assign rcache_line[6][41].status_reg.re    = reg2hw.status_1577.re;


  assign rcache_line[6][42].tag_reg.tag      = reg2hw.tag_1578.q;
  assign rcache_line[6][42].tag_reg.qe       = reg2hw.tag_1578.qe;
  assign rcache_line[6][42].tag_reg.re       = reg2hw.tag_1578.re;
  assign rcache_line[6][42].status_reg.status = reg2hw.status_1578.q;//status_reg_t'(reg2hw.status_1578.q);
  assign rcache_line[6][42].status_reg.qe    = reg2hw.status_1578.qe;
  assign rcache_line[6][42].status_reg.re    = reg2hw.status_1578.re;


  assign rcache_line[6][43].tag_reg.tag      = reg2hw.tag_1579.q;
  assign rcache_line[6][43].tag_reg.qe       = reg2hw.tag_1579.qe;
  assign rcache_line[6][43].tag_reg.re       = reg2hw.tag_1579.re;
  assign rcache_line[6][43].status_reg.status = reg2hw.status_1579.q;//status_reg_t'(reg2hw.status_1579.q);
  assign rcache_line[6][43].status_reg.qe    = reg2hw.status_1579.qe;
  assign rcache_line[6][43].status_reg.re    = reg2hw.status_1579.re;


  assign rcache_line[6][44].tag_reg.tag      = reg2hw.tag_1580.q;
  assign rcache_line[6][44].tag_reg.qe       = reg2hw.tag_1580.qe;
  assign rcache_line[6][44].tag_reg.re       = reg2hw.tag_1580.re;
  assign rcache_line[6][44].status_reg.status = reg2hw.status_1580.q;//status_reg_t'(reg2hw.status_1580.q);
  assign rcache_line[6][44].status_reg.qe    = reg2hw.status_1580.qe;
  assign rcache_line[6][44].status_reg.re    = reg2hw.status_1580.re;


  assign rcache_line[6][45].tag_reg.tag      = reg2hw.tag_1581.q;
  assign rcache_line[6][45].tag_reg.qe       = reg2hw.tag_1581.qe;
  assign rcache_line[6][45].tag_reg.re       = reg2hw.tag_1581.re;
  assign rcache_line[6][45].status_reg.status = reg2hw.status_1581.q;//status_reg_t'(reg2hw.status_1581.q);
  assign rcache_line[6][45].status_reg.qe    = reg2hw.status_1581.qe;
  assign rcache_line[6][45].status_reg.re    = reg2hw.status_1581.re;


  assign rcache_line[6][46].tag_reg.tag      = reg2hw.tag_1582.q;
  assign rcache_line[6][46].tag_reg.qe       = reg2hw.tag_1582.qe;
  assign rcache_line[6][46].tag_reg.re       = reg2hw.tag_1582.re;
  assign rcache_line[6][46].status_reg.status = reg2hw.status_1582.q;//status_reg_t'(reg2hw.status_1582.q);
  assign rcache_line[6][46].status_reg.qe    = reg2hw.status_1582.qe;
  assign rcache_line[6][46].status_reg.re    = reg2hw.status_1582.re;


  assign rcache_line[6][47].tag_reg.tag      = reg2hw.tag_1583.q;
  assign rcache_line[6][47].tag_reg.qe       = reg2hw.tag_1583.qe;
  assign rcache_line[6][47].tag_reg.re       = reg2hw.tag_1583.re;
  assign rcache_line[6][47].status_reg.status = reg2hw.status_1583.q;//status_reg_t'(reg2hw.status_1583.q);
  assign rcache_line[6][47].status_reg.qe    = reg2hw.status_1583.qe;
  assign rcache_line[6][47].status_reg.re    = reg2hw.status_1583.re;


  assign rcache_line[6][48].tag_reg.tag      = reg2hw.tag_1584.q;
  assign rcache_line[6][48].tag_reg.qe       = reg2hw.tag_1584.qe;
  assign rcache_line[6][48].tag_reg.re       = reg2hw.tag_1584.re;
  assign rcache_line[6][48].status_reg.status = reg2hw.status_1584.q;//status_reg_t'(reg2hw.status_1584.q);
  assign rcache_line[6][48].status_reg.qe    = reg2hw.status_1584.qe;
  assign rcache_line[6][48].status_reg.re    = reg2hw.status_1584.re;


  assign rcache_line[6][49].tag_reg.tag      = reg2hw.tag_1585.q;
  assign rcache_line[6][49].tag_reg.qe       = reg2hw.tag_1585.qe;
  assign rcache_line[6][49].tag_reg.re       = reg2hw.tag_1585.re;
  assign rcache_line[6][49].status_reg.status = reg2hw.status_1585.q;//status_reg_t'(reg2hw.status_1585.q);
  assign rcache_line[6][49].status_reg.qe    = reg2hw.status_1585.qe;
  assign rcache_line[6][49].status_reg.re    = reg2hw.status_1585.re;


  assign rcache_line[6][50].tag_reg.tag      = reg2hw.tag_1586.q;
  assign rcache_line[6][50].tag_reg.qe       = reg2hw.tag_1586.qe;
  assign rcache_line[6][50].tag_reg.re       = reg2hw.tag_1586.re;
  assign rcache_line[6][50].status_reg.status = reg2hw.status_1586.q;//status_reg_t'(reg2hw.status_1586.q);
  assign rcache_line[6][50].status_reg.qe    = reg2hw.status_1586.qe;
  assign rcache_line[6][50].status_reg.re    = reg2hw.status_1586.re;


  assign rcache_line[6][51].tag_reg.tag      = reg2hw.tag_1587.q;
  assign rcache_line[6][51].tag_reg.qe       = reg2hw.tag_1587.qe;
  assign rcache_line[6][51].tag_reg.re       = reg2hw.tag_1587.re;
  assign rcache_line[6][51].status_reg.status = reg2hw.status_1587.q;//status_reg_t'(reg2hw.status_1587.q);
  assign rcache_line[6][51].status_reg.qe    = reg2hw.status_1587.qe;
  assign rcache_line[6][51].status_reg.re    = reg2hw.status_1587.re;


  assign rcache_line[6][52].tag_reg.tag      = reg2hw.tag_1588.q;
  assign rcache_line[6][52].tag_reg.qe       = reg2hw.tag_1588.qe;
  assign rcache_line[6][52].tag_reg.re       = reg2hw.tag_1588.re;
  assign rcache_line[6][52].status_reg.status = reg2hw.status_1588.q;//status_reg_t'(reg2hw.status_1588.q);
  assign rcache_line[6][52].status_reg.qe    = reg2hw.status_1588.qe;
  assign rcache_line[6][52].status_reg.re    = reg2hw.status_1588.re;


  assign rcache_line[6][53].tag_reg.tag      = reg2hw.tag_1589.q;
  assign rcache_line[6][53].tag_reg.qe       = reg2hw.tag_1589.qe;
  assign rcache_line[6][53].tag_reg.re       = reg2hw.tag_1589.re;
  assign rcache_line[6][53].status_reg.status = reg2hw.status_1589.q;//status_reg_t'(reg2hw.status_1589.q);
  assign rcache_line[6][53].status_reg.qe    = reg2hw.status_1589.qe;
  assign rcache_line[6][53].status_reg.re    = reg2hw.status_1589.re;


  assign rcache_line[6][54].tag_reg.tag      = reg2hw.tag_1590.q;
  assign rcache_line[6][54].tag_reg.qe       = reg2hw.tag_1590.qe;
  assign rcache_line[6][54].tag_reg.re       = reg2hw.tag_1590.re;
  assign rcache_line[6][54].status_reg.status = reg2hw.status_1590.q;//status_reg_t'(reg2hw.status_1590.q);
  assign rcache_line[6][54].status_reg.qe    = reg2hw.status_1590.qe;
  assign rcache_line[6][54].status_reg.re    = reg2hw.status_1590.re;


  assign rcache_line[6][55].tag_reg.tag      = reg2hw.tag_1591.q;
  assign rcache_line[6][55].tag_reg.qe       = reg2hw.tag_1591.qe;
  assign rcache_line[6][55].tag_reg.re       = reg2hw.tag_1591.re;
  assign rcache_line[6][55].status_reg.status = reg2hw.status_1591.q;//status_reg_t'(reg2hw.status_1591.q);
  assign rcache_line[6][55].status_reg.qe    = reg2hw.status_1591.qe;
  assign rcache_line[6][55].status_reg.re    = reg2hw.status_1591.re;


  assign rcache_line[6][56].tag_reg.tag      = reg2hw.tag_1592.q;
  assign rcache_line[6][56].tag_reg.qe       = reg2hw.tag_1592.qe;
  assign rcache_line[6][56].tag_reg.re       = reg2hw.tag_1592.re;
  assign rcache_line[6][56].status_reg.status = reg2hw.status_1592.q;//status_reg_t'(reg2hw.status_1592.q);
  assign rcache_line[6][56].status_reg.qe    = reg2hw.status_1592.qe;
  assign rcache_line[6][56].status_reg.re    = reg2hw.status_1592.re;


  assign rcache_line[6][57].tag_reg.tag      = reg2hw.tag_1593.q;
  assign rcache_line[6][57].tag_reg.qe       = reg2hw.tag_1593.qe;
  assign rcache_line[6][57].tag_reg.re       = reg2hw.tag_1593.re;
  assign rcache_line[6][57].status_reg.status = reg2hw.status_1593.q;//status_reg_t'(reg2hw.status_1593.q);
  assign rcache_line[6][57].status_reg.qe    = reg2hw.status_1593.qe;
  assign rcache_line[6][57].status_reg.re    = reg2hw.status_1593.re;


  assign rcache_line[6][58].tag_reg.tag      = reg2hw.tag_1594.q;
  assign rcache_line[6][58].tag_reg.qe       = reg2hw.tag_1594.qe;
  assign rcache_line[6][58].tag_reg.re       = reg2hw.tag_1594.re;
  assign rcache_line[6][58].status_reg.status = reg2hw.status_1594.q;//status_reg_t'(reg2hw.status_1594.q);
  assign rcache_line[6][58].status_reg.qe    = reg2hw.status_1594.qe;
  assign rcache_line[6][58].status_reg.re    = reg2hw.status_1594.re;


  assign rcache_line[6][59].tag_reg.tag      = reg2hw.tag_1595.q;
  assign rcache_line[6][59].tag_reg.qe       = reg2hw.tag_1595.qe;
  assign rcache_line[6][59].tag_reg.re       = reg2hw.tag_1595.re;
  assign rcache_line[6][59].status_reg.status = reg2hw.status_1595.q;//status_reg_t'(reg2hw.status_1595.q);
  assign rcache_line[6][59].status_reg.qe    = reg2hw.status_1595.qe;
  assign rcache_line[6][59].status_reg.re    = reg2hw.status_1595.re;


  assign rcache_line[6][60].tag_reg.tag      = reg2hw.tag_1596.q;
  assign rcache_line[6][60].tag_reg.qe       = reg2hw.tag_1596.qe;
  assign rcache_line[6][60].tag_reg.re       = reg2hw.tag_1596.re;
  assign rcache_line[6][60].status_reg.status = reg2hw.status_1596.q;//status_reg_t'(reg2hw.status_1596.q);
  assign rcache_line[6][60].status_reg.qe    = reg2hw.status_1596.qe;
  assign rcache_line[6][60].status_reg.re    = reg2hw.status_1596.re;


  assign rcache_line[6][61].tag_reg.tag      = reg2hw.tag_1597.q;
  assign rcache_line[6][61].tag_reg.qe       = reg2hw.tag_1597.qe;
  assign rcache_line[6][61].tag_reg.re       = reg2hw.tag_1597.re;
  assign rcache_line[6][61].status_reg.status = reg2hw.status_1597.q;//status_reg_t'(reg2hw.status_1597.q);
  assign rcache_line[6][61].status_reg.qe    = reg2hw.status_1597.qe;
  assign rcache_line[6][61].status_reg.re    = reg2hw.status_1597.re;


  assign rcache_line[6][62].tag_reg.tag      = reg2hw.tag_1598.q;
  assign rcache_line[6][62].tag_reg.qe       = reg2hw.tag_1598.qe;
  assign rcache_line[6][62].tag_reg.re       = reg2hw.tag_1598.re;
  assign rcache_line[6][62].status_reg.status = reg2hw.status_1598.q;//status_reg_t'(reg2hw.status_1598.q);
  assign rcache_line[6][62].status_reg.qe    = reg2hw.status_1598.qe;
  assign rcache_line[6][62].status_reg.re    = reg2hw.status_1598.re;


  assign rcache_line[6][63].tag_reg.tag      = reg2hw.tag_1599.q;
  assign rcache_line[6][63].tag_reg.qe       = reg2hw.tag_1599.qe;
  assign rcache_line[6][63].tag_reg.re       = reg2hw.tag_1599.re;
  assign rcache_line[6][63].status_reg.status = reg2hw.status_1599.q;//status_reg_t'(reg2hw.status_1599.q);
  assign rcache_line[6][63].status_reg.qe    = reg2hw.status_1599.qe;
  assign rcache_line[6][63].status_reg.re    = reg2hw.status_1599.re;


  assign rcache_line[6][64].tag_reg.tag      = reg2hw.tag_1600.q;
  assign rcache_line[6][64].tag_reg.qe       = reg2hw.tag_1600.qe;
  assign rcache_line[6][64].tag_reg.re       = reg2hw.tag_1600.re;
  assign rcache_line[6][64].status_reg.status = reg2hw.status_1600.q;//status_reg_t'(reg2hw.status_1600.q);
  assign rcache_line[6][64].status_reg.qe    = reg2hw.status_1600.qe;
  assign rcache_line[6][64].status_reg.re    = reg2hw.status_1600.re;


  assign rcache_line[6][65].tag_reg.tag      = reg2hw.tag_1601.q;
  assign rcache_line[6][65].tag_reg.qe       = reg2hw.tag_1601.qe;
  assign rcache_line[6][65].tag_reg.re       = reg2hw.tag_1601.re;
  assign rcache_line[6][65].status_reg.status = reg2hw.status_1601.q;//status_reg_t'(reg2hw.status_1601.q);
  assign rcache_line[6][65].status_reg.qe    = reg2hw.status_1601.qe;
  assign rcache_line[6][65].status_reg.re    = reg2hw.status_1601.re;


  assign rcache_line[6][66].tag_reg.tag      = reg2hw.tag_1602.q;
  assign rcache_line[6][66].tag_reg.qe       = reg2hw.tag_1602.qe;
  assign rcache_line[6][66].tag_reg.re       = reg2hw.tag_1602.re;
  assign rcache_line[6][66].status_reg.status = reg2hw.status_1602.q;//status_reg_t'(reg2hw.status_1602.q);
  assign rcache_line[6][66].status_reg.qe    = reg2hw.status_1602.qe;
  assign rcache_line[6][66].status_reg.re    = reg2hw.status_1602.re;


  assign rcache_line[6][67].tag_reg.tag      = reg2hw.tag_1603.q;
  assign rcache_line[6][67].tag_reg.qe       = reg2hw.tag_1603.qe;
  assign rcache_line[6][67].tag_reg.re       = reg2hw.tag_1603.re;
  assign rcache_line[6][67].status_reg.status = reg2hw.status_1603.q;//status_reg_t'(reg2hw.status_1603.q);
  assign rcache_line[6][67].status_reg.qe    = reg2hw.status_1603.qe;
  assign rcache_line[6][67].status_reg.re    = reg2hw.status_1603.re;


  assign rcache_line[6][68].tag_reg.tag      = reg2hw.tag_1604.q;
  assign rcache_line[6][68].tag_reg.qe       = reg2hw.tag_1604.qe;
  assign rcache_line[6][68].tag_reg.re       = reg2hw.tag_1604.re;
  assign rcache_line[6][68].status_reg.status = reg2hw.status_1604.q;//status_reg_t'(reg2hw.status_1604.q);
  assign rcache_line[6][68].status_reg.qe    = reg2hw.status_1604.qe;
  assign rcache_line[6][68].status_reg.re    = reg2hw.status_1604.re;


  assign rcache_line[6][69].tag_reg.tag      = reg2hw.tag_1605.q;
  assign rcache_line[6][69].tag_reg.qe       = reg2hw.tag_1605.qe;
  assign rcache_line[6][69].tag_reg.re       = reg2hw.tag_1605.re;
  assign rcache_line[6][69].status_reg.status = reg2hw.status_1605.q;//status_reg_t'(reg2hw.status_1605.q);
  assign rcache_line[6][69].status_reg.qe    = reg2hw.status_1605.qe;
  assign rcache_line[6][69].status_reg.re    = reg2hw.status_1605.re;


  assign rcache_line[6][70].tag_reg.tag      = reg2hw.tag_1606.q;
  assign rcache_line[6][70].tag_reg.qe       = reg2hw.tag_1606.qe;
  assign rcache_line[6][70].tag_reg.re       = reg2hw.tag_1606.re;
  assign rcache_line[6][70].status_reg.status = reg2hw.status_1606.q;//status_reg_t'(reg2hw.status_1606.q);
  assign rcache_line[6][70].status_reg.qe    = reg2hw.status_1606.qe;
  assign rcache_line[6][70].status_reg.re    = reg2hw.status_1606.re;


  assign rcache_line[6][71].tag_reg.tag      = reg2hw.tag_1607.q;
  assign rcache_line[6][71].tag_reg.qe       = reg2hw.tag_1607.qe;
  assign rcache_line[6][71].tag_reg.re       = reg2hw.tag_1607.re;
  assign rcache_line[6][71].status_reg.status = reg2hw.status_1607.q;//status_reg_t'(reg2hw.status_1607.q);
  assign rcache_line[6][71].status_reg.qe    = reg2hw.status_1607.qe;
  assign rcache_line[6][71].status_reg.re    = reg2hw.status_1607.re;


  assign rcache_line[6][72].tag_reg.tag      = reg2hw.tag_1608.q;
  assign rcache_line[6][72].tag_reg.qe       = reg2hw.tag_1608.qe;
  assign rcache_line[6][72].tag_reg.re       = reg2hw.tag_1608.re;
  assign rcache_line[6][72].status_reg.status = reg2hw.status_1608.q;//status_reg_t'(reg2hw.status_1608.q);
  assign rcache_line[6][72].status_reg.qe    = reg2hw.status_1608.qe;
  assign rcache_line[6][72].status_reg.re    = reg2hw.status_1608.re;


  assign rcache_line[6][73].tag_reg.tag      = reg2hw.tag_1609.q;
  assign rcache_line[6][73].tag_reg.qe       = reg2hw.tag_1609.qe;
  assign rcache_line[6][73].tag_reg.re       = reg2hw.tag_1609.re;
  assign rcache_line[6][73].status_reg.status = reg2hw.status_1609.q;//status_reg_t'(reg2hw.status_1609.q);
  assign rcache_line[6][73].status_reg.qe    = reg2hw.status_1609.qe;
  assign rcache_line[6][73].status_reg.re    = reg2hw.status_1609.re;


  assign rcache_line[6][74].tag_reg.tag      = reg2hw.tag_1610.q;
  assign rcache_line[6][74].tag_reg.qe       = reg2hw.tag_1610.qe;
  assign rcache_line[6][74].tag_reg.re       = reg2hw.tag_1610.re;
  assign rcache_line[6][74].status_reg.status = reg2hw.status_1610.q;//status_reg_t'(reg2hw.status_1610.q);
  assign rcache_line[6][74].status_reg.qe    = reg2hw.status_1610.qe;
  assign rcache_line[6][74].status_reg.re    = reg2hw.status_1610.re;


  assign rcache_line[6][75].tag_reg.tag      = reg2hw.tag_1611.q;
  assign rcache_line[6][75].tag_reg.qe       = reg2hw.tag_1611.qe;
  assign rcache_line[6][75].tag_reg.re       = reg2hw.tag_1611.re;
  assign rcache_line[6][75].status_reg.status = reg2hw.status_1611.q;//status_reg_t'(reg2hw.status_1611.q);
  assign rcache_line[6][75].status_reg.qe    = reg2hw.status_1611.qe;
  assign rcache_line[6][75].status_reg.re    = reg2hw.status_1611.re;


  assign rcache_line[6][76].tag_reg.tag      = reg2hw.tag_1612.q;
  assign rcache_line[6][76].tag_reg.qe       = reg2hw.tag_1612.qe;
  assign rcache_line[6][76].tag_reg.re       = reg2hw.tag_1612.re;
  assign rcache_line[6][76].status_reg.status = reg2hw.status_1612.q;//status_reg_t'(reg2hw.status_1612.q);
  assign rcache_line[6][76].status_reg.qe    = reg2hw.status_1612.qe;
  assign rcache_line[6][76].status_reg.re    = reg2hw.status_1612.re;


  assign rcache_line[6][77].tag_reg.tag      = reg2hw.tag_1613.q;
  assign rcache_line[6][77].tag_reg.qe       = reg2hw.tag_1613.qe;
  assign rcache_line[6][77].tag_reg.re       = reg2hw.tag_1613.re;
  assign rcache_line[6][77].status_reg.status = reg2hw.status_1613.q;//status_reg_t'(reg2hw.status_1613.q);
  assign rcache_line[6][77].status_reg.qe    = reg2hw.status_1613.qe;
  assign rcache_line[6][77].status_reg.re    = reg2hw.status_1613.re;


  assign rcache_line[6][78].tag_reg.tag      = reg2hw.tag_1614.q;
  assign rcache_line[6][78].tag_reg.qe       = reg2hw.tag_1614.qe;
  assign rcache_line[6][78].tag_reg.re       = reg2hw.tag_1614.re;
  assign rcache_line[6][78].status_reg.status = reg2hw.status_1614.q;//status_reg_t'(reg2hw.status_1614.q);
  assign rcache_line[6][78].status_reg.qe    = reg2hw.status_1614.qe;
  assign rcache_line[6][78].status_reg.re    = reg2hw.status_1614.re;


  assign rcache_line[6][79].tag_reg.tag      = reg2hw.tag_1615.q;
  assign rcache_line[6][79].tag_reg.qe       = reg2hw.tag_1615.qe;
  assign rcache_line[6][79].tag_reg.re       = reg2hw.tag_1615.re;
  assign rcache_line[6][79].status_reg.status = reg2hw.status_1615.q;//status_reg_t'(reg2hw.status_1615.q);
  assign rcache_line[6][79].status_reg.qe    = reg2hw.status_1615.qe;
  assign rcache_line[6][79].status_reg.re    = reg2hw.status_1615.re;


  assign rcache_line[6][80].tag_reg.tag      = reg2hw.tag_1616.q;
  assign rcache_line[6][80].tag_reg.qe       = reg2hw.tag_1616.qe;
  assign rcache_line[6][80].tag_reg.re       = reg2hw.tag_1616.re;
  assign rcache_line[6][80].status_reg.status = reg2hw.status_1616.q;//status_reg_t'(reg2hw.status_1616.q);
  assign rcache_line[6][80].status_reg.qe    = reg2hw.status_1616.qe;
  assign rcache_line[6][80].status_reg.re    = reg2hw.status_1616.re;


  assign rcache_line[6][81].tag_reg.tag      = reg2hw.tag_1617.q;
  assign rcache_line[6][81].tag_reg.qe       = reg2hw.tag_1617.qe;
  assign rcache_line[6][81].tag_reg.re       = reg2hw.tag_1617.re;
  assign rcache_line[6][81].status_reg.status = reg2hw.status_1617.q;//status_reg_t'(reg2hw.status_1617.q);
  assign rcache_line[6][81].status_reg.qe    = reg2hw.status_1617.qe;
  assign rcache_line[6][81].status_reg.re    = reg2hw.status_1617.re;


  assign rcache_line[6][82].tag_reg.tag      = reg2hw.tag_1618.q;
  assign rcache_line[6][82].tag_reg.qe       = reg2hw.tag_1618.qe;
  assign rcache_line[6][82].tag_reg.re       = reg2hw.tag_1618.re;
  assign rcache_line[6][82].status_reg.status = reg2hw.status_1618.q;//status_reg_t'(reg2hw.status_1618.q);
  assign rcache_line[6][82].status_reg.qe    = reg2hw.status_1618.qe;
  assign rcache_line[6][82].status_reg.re    = reg2hw.status_1618.re;


  assign rcache_line[6][83].tag_reg.tag      = reg2hw.tag_1619.q;
  assign rcache_line[6][83].tag_reg.qe       = reg2hw.tag_1619.qe;
  assign rcache_line[6][83].tag_reg.re       = reg2hw.tag_1619.re;
  assign rcache_line[6][83].status_reg.status = reg2hw.status_1619.q;//status_reg_t'(reg2hw.status_1619.q);
  assign rcache_line[6][83].status_reg.qe    = reg2hw.status_1619.qe;
  assign rcache_line[6][83].status_reg.re    = reg2hw.status_1619.re;


  assign rcache_line[6][84].tag_reg.tag      = reg2hw.tag_1620.q;
  assign rcache_line[6][84].tag_reg.qe       = reg2hw.tag_1620.qe;
  assign rcache_line[6][84].tag_reg.re       = reg2hw.tag_1620.re;
  assign rcache_line[6][84].status_reg.status = reg2hw.status_1620.q;//status_reg_t'(reg2hw.status_1620.q);
  assign rcache_line[6][84].status_reg.qe    = reg2hw.status_1620.qe;
  assign rcache_line[6][84].status_reg.re    = reg2hw.status_1620.re;


  assign rcache_line[6][85].tag_reg.tag      = reg2hw.tag_1621.q;
  assign rcache_line[6][85].tag_reg.qe       = reg2hw.tag_1621.qe;
  assign rcache_line[6][85].tag_reg.re       = reg2hw.tag_1621.re;
  assign rcache_line[6][85].status_reg.status = reg2hw.status_1621.q;//status_reg_t'(reg2hw.status_1621.q);
  assign rcache_line[6][85].status_reg.qe    = reg2hw.status_1621.qe;
  assign rcache_line[6][85].status_reg.re    = reg2hw.status_1621.re;


  assign rcache_line[6][86].tag_reg.tag      = reg2hw.tag_1622.q;
  assign rcache_line[6][86].tag_reg.qe       = reg2hw.tag_1622.qe;
  assign rcache_line[6][86].tag_reg.re       = reg2hw.tag_1622.re;
  assign rcache_line[6][86].status_reg.status = reg2hw.status_1622.q;//status_reg_t'(reg2hw.status_1622.q);
  assign rcache_line[6][86].status_reg.qe    = reg2hw.status_1622.qe;
  assign rcache_line[6][86].status_reg.re    = reg2hw.status_1622.re;


  assign rcache_line[6][87].tag_reg.tag      = reg2hw.tag_1623.q;
  assign rcache_line[6][87].tag_reg.qe       = reg2hw.tag_1623.qe;
  assign rcache_line[6][87].tag_reg.re       = reg2hw.tag_1623.re;
  assign rcache_line[6][87].status_reg.status = reg2hw.status_1623.q;//status_reg_t'(reg2hw.status_1623.q);
  assign rcache_line[6][87].status_reg.qe    = reg2hw.status_1623.qe;
  assign rcache_line[6][87].status_reg.re    = reg2hw.status_1623.re;


  assign rcache_line[6][88].tag_reg.tag      = reg2hw.tag_1624.q;
  assign rcache_line[6][88].tag_reg.qe       = reg2hw.tag_1624.qe;
  assign rcache_line[6][88].tag_reg.re       = reg2hw.tag_1624.re;
  assign rcache_line[6][88].status_reg.status = reg2hw.status_1624.q;//status_reg_t'(reg2hw.status_1624.q);
  assign rcache_line[6][88].status_reg.qe    = reg2hw.status_1624.qe;
  assign rcache_line[6][88].status_reg.re    = reg2hw.status_1624.re;


  assign rcache_line[6][89].tag_reg.tag      = reg2hw.tag_1625.q;
  assign rcache_line[6][89].tag_reg.qe       = reg2hw.tag_1625.qe;
  assign rcache_line[6][89].tag_reg.re       = reg2hw.tag_1625.re;
  assign rcache_line[6][89].status_reg.status = reg2hw.status_1625.q;//status_reg_t'(reg2hw.status_1625.q);
  assign rcache_line[6][89].status_reg.qe    = reg2hw.status_1625.qe;
  assign rcache_line[6][89].status_reg.re    = reg2hw.status_1625.re;


  assign rcache_line[6][90].tag_reg.tag      = reg2hw.tag_1626.q;
  assign rcache_line[6][90].tag_reg.qe       = reg2hw.tag_1626.qe;
  assign rcache_line[6][90].tag_reg.re       = reg2hw.tag_1626.re;
  assign rcache_line[6][90].status_reg.status = reg2hw.status_1626.q;//status_reg_t'(reg2hw.status_1626.q);
  assign rcache_line[6][90].status_reg.qe    = reg2hw.status_1626.qe;
  assign rcache_line[6][90].status_reg.re    = reg2hw.status_1626.re;


  assign rcache_line[6][91].tag_reg.tag      = reg2hw.tag_1627.q;
  assign rcache_line[6][91].tag_reg.qe       = reg2hw.tag_1627.qe;
  assign rcache_line[6][91].tag_reg.re       = reg2hw.tag_1627.re;
  assign rcache_line[6][91].status_reg.status = reg2hw.status_1627.q;//status_reg_t'(reg2hw.status_1627.q);
  assign rcache_line[6][91].status_reg.qe    = reg2hw.status_1627.qe;
  assign rcache_line[6][91].status_reg.re    = reg2hw.status_1627.re;


  assign rcache_line[6][92].tag_reg.tag      = reg2hw.tag_1628.q;
  assign rcache_line[6][92].tag_reg.qe       = reg2hw.tag_1628.qe;
  assign rcache_line[6][92].tag_reg.re       = reg2hw.tag_1628.re;
  assign rcache_line[6][92].status_reg.status = reg2hw.status_1628.q;//status_reg_t'(reg2hw.status_1628.q);
  assign rcache_line[6][92].status_reg.qe    = reg2hw.status_1628.qe;
  assign rcache_line[6][92].status_reg.re    = reg2hw.status_1628.re;


  assign rcache_line[6][93].tag_reg.tag      = reg2hw.tag_1629.q;
  assign rcache_line[6][93].tag_reg.qe       = reg2hw.tag_1629.qe;
  assign rcache_line[6][93].tag_reg.re       = reg2hw.tag_1629.re;
  assign rcache_line[6][93].status_reg.status = reg2hw.status_1629.q;//status_reg_t'(reg2hw.status_1629.q);
  assign rcache_line[6][93].status_reg.qe    = reg2hw.status_1629.qe;
  assign rcache_line[6][93].status_reg.re    = reg2hw.status_1629.re;


  assign rcache_line[6][94].tag_reg.tag      = reg2hw.tag_1630.q;
  assign rcache_line[6][94].tag_reg.qe       = reg2hw.tag_1630.qe;
  assign rcache_line[6][94].tag_reg.re       = reg2hw.tag_1630.re;
  assign rcache_line[6][94].status_reg.status = reg2hw.status_1630.q;//status_reg_t'(reg2hw.status_1630.q);
  assign rcache_line[6][94].status_reg.qe    = reg2hw.status_1630.qe;
  assign rcache_line[6][94].status_reg.re    = reg2hw.status_1630.re;


  assign rcache_line[6][95].tag_reg.tag      = reg2hw.tag_1631.q;
  assign rcache_line[6][95].tag_reg.qe       = reg2hw.tag_1631.qe;
  assign rcache_line[6][95].tag_reg.re       = reg2hw.tag_1631.re;
  assign rcache_line[6][95].status_reg.status = reg2hw.status_1631.q;//status_reg_t'(reg2hw.status_1631.q);
  assign rcache_line[6][95].status_reg.qe    = reg2hw.status_1631.qe;
  assign rcache_line[6][95].status_reg.re    = reg2hw.status_1631.re;


  assign rcache_line[6][96].tag_reg.tag      = reg2hw.tag_1632.q;
  assign rcache_line[6][96].tag_reg.qe       = reg2hw.tag_1632.qe;
  assign rcache_line[6][96].tag_reg.re       = reg2hw.tag_1632.re;
  assign rcache_line[6][96].status_reg.status = reg2hw.status_1632.q;//status_reg_t'(reg2hw.status_1632.q);
  assign rcache_line[6][96].status_reg.qe    = reg2hw.status_1632.qe;
  assign rcache_line[6][96].status_reg.re    = reg2hw.status_1632.re;


  assign rcache_line[6][97].tag_reg.tag      = reg2hw.tag_1633.q;
  assign rcache_line[6][97].tag_reg.qe       = reg2hw.tag_1633.qe;
  assign rcache_line[6][97].tag_reg.re       = reg2hw.tag_1633.re;
  assign rcache_line[6][97].status_reg.status = reg2hw.status_1633.q;//status_reg_t'(reg2hw.status_1633.q);
  assign rcache_line[6][97].status_reg.qe    = reg2hw.status_1633.qe;
  assign rcache_line[6][97].status_reg.re    = reg2hw.status_1633.re;


  assign rcache_line[6][98].tag_reg.tag      = reg2hw.tag_1634.q;
  assign rcache_line[6][98].tag_reg.qe       = reg2hw.tag_1634.qe;
  assign rcache_line[6][98].tag_reg.re       = reg2hw.tag_1634.re;
  assign rcache_line[6][98].status_reg.status = reg2hw.status_1634.q;//status_reg_t'(reg2hw.status_1634.q);
  assign rcache_line[6][98].status_reg.qe    = reg2hw.status_1634.qe;
  assign rcache_line[6][98].status_reg.re    = reg2hw.status_1634.re;


  assign rcache_line[6][99].tag_reg.tag      = reg2hw.tag_1635.q;
  assign rcache_line[6][99].tag_reg.qe       = reg2hw.tag_1635.qe;
  assign rcache_line[6][99].tag_reg.re       = reg2hw.tag_1635.re;
  assign rcache_line[6][99].status_reg.status = reg2hw.status_1635.q;//status_reg_t'(reg2hw.status_1635.q);
  assign rcache_line[6][99].status_reg.qe    = reg2hw.status_1635.qe;
  assign rcache_line[6][99].status_reg.re    = reg2hw.status_1635.re;


  assign rcache_line[6][100].tag_reg.tag      = reg2hw.tag_1636.q;
  assign rcache_line[6][100].tag_reg.qe       = reg2hw.tag_1636.qe;
  assign rcache_line[6][100].tag_reg.re       = reg2hw.tag_1636.re;
  assign rcache_line[6][100].status_reg.status = reg2hw.status_1636.q;//status_reg_t'(reg2hw.status_1636.q);
  assign rcache_line[6][100].status_reg.qe    = reg2hw.status_1636.qe;
  assign rcache_line[6][100].status_reg.re    = reg2hw.status_1636.re;


  assign rcache_line[6][101].tag_reg.tag      = reg2hw.tag_1637.q;
  assign rcache_line[6][101].tag_reg.qe       = reg2hw.tag_1637.qe;
  assign rcache_line[6][101].tag_reg.re       = reg2hw.tag_1637.re;
  assign rcache_line[6][101].status_reg.status = reg2hw.status_1637.q;//status_reg_t'(reg2hw.status_1637.q);
  assign rcache_line[6][101].status_reg.qe    = reg2hw.status_1637.qe;
  assign rcache_line[6][101].status_reg.re    = reg2hw.status_1637.re;


  assign rcache_line[6][102].tag_reg.tag      = reg2hw.tag_1638.q;
  assign rcache_line[6][102].tag_reg.qe       = reg2hw.tag_1638.qe;
  assign rcache_line[6][102].tag_reg.re       = reg2hw.tag_1638.re;
  assign rcache_line[6][102].status_reg.status = reg2hw.status_1638.q;//status_reg_t'(reg2hw.status_1638.q);
  assign rcache_line[6][102].status_reg.qe    = reg2hw.status_1638.qe;
  assign rcache_line[6][102].status_reg.re    = reg2hw.status_1638.re;


  assign rcache_line[6][103].tag_reg.tag      = reg2hw.tag_1639.q;
  assign rcache_line[6][103].tag_reg.qe       = reg2hw.tag_1639.qe;
  assign rcache_line[6][103].tag_reg.re       = reg2hw.tag_1639.re;
  assign rcache_line[6][103].status_reg.status = reg2hw.status_1639.q;//status_reg_t'(reg2hw.status_1639.q);
  assign rcache_line[6][103].status_reg.qe    = reg2hw.status_1639.qe;
  assign rcache_line[6][103].status_reg.re    = reg2hw.status_1639.re;


  assign rcache_line[6][104].tag_reg.tag      = reg2hw.tag_1640.q;
  assign rcache_line[6][104].tag_reg.qe       = reg2hw.tag_1640.qe;
  assign rcache_line[6][104].tag_reg.re       = reg2hw.tag_1640.re;
  assign rcache_line[6][104].status_reg.status = reg2hw.status_1640.q;//status_reg_t'(reg2hw.status_1640.q);
  assign rcache_line[6][104].status_reg.qe    = reg2hw.status_1640.qe;
  assign rcache_line[6][104].status_reg.re    = reg2hw.status_1640.re;


  assign rcache_line[6][105].tag_reg.tag      = reg2hw.tag_1641.q;
  assign rcache_line[6][105].tag_reg.qe       = reg2hw.tag_1641.qe;
  assign rcache_line[6][105].tag_reg.re       = reg2hw.tag_1641.re;
  assign rcache_line[6][105].status_reg.status = reg2hw.status_1641.q;//status_reg_t'(reg2hw.status_1641.q);
  assign rcache_line[6][105].status_reg.qe    = reg2hw.status_1641.qe;
  assign rcache_line[6][105].status_reg.re    = reg2hw.status_1641.re;


  assign rcache_line[6][106].tag_reg.tag      = reg2hw.tag_1642.q;
  assign rcache_line[6][106].tag_reg.qe       = reg2hw.tag_1642.qe;
  assign rcache_line[6][106].tag_reg.re       = reg2hw.tag_1642.re;
  assign rcache_line[6][106].status_reg.status = reg2hw.status_1642.q;//status_reg_t'(reg2hw.status_1642.q);
  assign rcache_line[6][106].status_reg.qe    = reg2hw.status_1642.qe;
  assign rcache_line[6][106].status_reg.re    = reg2hw.status_1642.re;


  assign rcache_line[6][107].tag_reg.tag      = reg2hw.tag_1643.q;
  assign rcache_line[6][107].tag_reg.qe       = reg2hw.tag_1643.qe;
  assign rcache_line[6][107].tag_reg.re       = reg2hw.tag_1643.re;
  assign rcache_line[6][107].status_reg.status = reg2hw.status_1643.q;//status_reg_t'(reg2hw.status_1643.q);
  assign rcache_line[6][107].status_reg.qe    = reg2hw.status_1643.qe;
  assign rcache_line[6][107].status_reg.re    = reg2hw.status_1643.re;


  assign rcache_line[6][108].tag_reg.tag      = reg2hw.tag_1644.q;
  assign rcache_line[6][108].tag_reg.qe       = reg2hw.tag_1644.qe;
  assign rcache_line[6][108].tag_reg.re       = reg2hw.tag_1644.re;
  assign rcache_line[6][108].status_reg.status = reg2hw.status_1644.q;//status_reg_t'(reg2hw.status_1644.q);
  assign rcache_line[6][108].status_reg.qe    = reg2hw.status_1644.qe;
  assign rcache_line[6][108].status_reg.re    = reg2hw.status_1644.re;


  assign rcache_line[6][109].tag_reg.tag      = reg2hw.tag_1645.q;
  assign rcache_line[6][109].tag_reg.qe       = reg2hw.tag_1645.qe;
  assign rcache_line[6][109].tag_reg.re       = reg2hw.tag_1645.re;
  assign rcache_line[6][109].status_reg.status = reg2hw.status_1645.q;//status_reg_t'(reg2hw.status_1645.q);
  assign rcache_line[6][109].status_reg.qe    = reg2hw.status_1645.qe;
  assign rcache_line[6][109].status_reg.re    = reg2hw.status_1645.re;


  assign rcache_line[6][110].tag_reg.tag      = reg2hw.tag_1646.q;
  assign rcache_line[6][110].tag_reg.qe       = reg2hw.tag_1646.qe;
  assign rcache_line[6][110].tag_reg.re       = reg2hw.tag_1646.re;
  assign rcache_line[6][110].status_reg.status = reg2hw.status_1646.q;//status_reg_t'(reg2hw.status_1646.q);
  assign rcache_line[6][110].status_reg.qe    = reg2hw.status_1646.qe;
  assign rcache_line[6][110].status_reg.re    = reg2hw.status_1646.re;


  assign rcache_line[6][111].tag_reg.tag      = reg2hw.tag_1647.q;
  assign rcache_line[6][111].tag_reg.qe       = reg2hw.tag_1647.qe;
  assign rcache_line[6][111].tag_reg.re       = reg2hw.tag_1647.re;
  assign rcache_line[6][111].status_reg.status = reg2hw.status_1647.q;//status_reg_t'(reg2hw.status_1647.q);
  assign rcache_line[6][111].status_reg.qe    = reg2hw.status_1647.qe;
  assign rcache_line[6][111].status_reg.re    = reg2hw.status_1647.re;


  assign rcache_line[6][112].tag_reg.tag      = reg2hw.tag_1648.q;
  assign rcache_line[6][112].tag_reg.qe       = reg2hw.tag_1648.qe;
  assign rcache_line[6][112].tag_reg.re       = reg2hw.tag_1648.re;
  assign rcache_line[6][112].status_reg.status = reg2hw.status_1648.q;//status_reg_t'(reg2hw.status_1648.q);
  assign rcache_line[6][112].status_reg.qe    = reg2hw.status_1648.qe;
  assign rcache_line[6][112].status_reg.re    = reg2hw.status_1648.re;


  assign rcache_line[6][113].tag_reg.tag      = reg2hw.tag_1649.q;
  assign rcache_line[6][113].tag_reg.qe       = reg2hw.tag_1649.qe;
  assign rcache_line[6][113].tag_reg.re       = reg2hw.tag_1649.re;
  assign rcache_line[6][113].status_reg.status = reg2hw.status_1649.q;//status_reg_t'(reg2hw.status_1649.q);
  assign rcache_line[6][113].status_reg.qe    = reg2hw.status_1649.qe;
  assign rcache_line[6][113].status_reg.re    = reg2hw.status_1649.re;


  assign rcache_line[6][114].tag_reg.tag      = reg2hw.tag_1650.q;
  assign rcache_line[6][114].tag_reg.qe       = reg2hw.tag_1650.qe;
  assign rcache_line[6][114].tag_reg.re       = reg2hw.tag_1650.re;
  assign rcache_line[6][114].status_reg.status = reg2hw.status_1650.q;//status_reg_t'(reg2hw.status_1650.q);
  assign rcache_line[6][114].status_reg.qe    = reg2hw.status_1650.qe;
  assign rcache_line[6][114].status_reg.re    = reg2hw.status_1650.re;


  assign rcache_line[6][115].tag_reg.tag      = reg2hw.tag_1651.q;
  assign rcache_line[6][115].tag_reg.qe       = reg2hw.tag_1651.qe;
  assign rcache_line[6][115].tag_reg.re       = reg2hw.tag_1651.re;
  assign rcache_line[6][115].status_reg.status = reg2hw.status_1651.q;//status_reg_t'(reg2hw.status_1651.q);
  assign rcache_line[6][115].status_reg.qe    = reg2hw.status_1651.qe;
  assign rcache_line[6][115].status_reg.re    = reg2hw.status_1651.re;


  assign rcache_line[6][116].tag_reg.tag      = reg2hw.tag_1652.q;
  assign rcache_line[6][116].tag_reg.qe       = reg2hw.tag_1652.qe;
  assign rcache_line[6][116].tag_reg.re       = reg2hw.tag_1652.re;
  assign rcache_line[6][116].status_reg.status = reg2hw.status_1652.q;//status_reg_t'(reg2hw.status_1652.q);
  assign rcache_line[6][116].status_reg.qe    = reg2hw.status_1652.qe;
  assign rcache_line[6][116].status_reg.re    = reg2hw.status_1652.re;


  assign rcache_line[6][117].tag_reg.tag      = reg2hw.tag_1653.q;
  assign rcache_line[6][117].tag_reg.qe       = reg2hw.tag_1653.qe;
  assign rcache_line[6][117].tag_reg.re       = reg2hw.tag_1653.re;
  assign rcache_line[6][117].status_reg.status = reg2hw.status_1653.q;//status_reg_t'(reg2hw.status_1653.q);
  assign rcache_line[6][117].status_reg.qe    = reg2hw.status_1653.qe;
  assign rcache_line[6][117].status_reg.re    = reg2hw.status_1653.re;


  assign rcache_line[6][118].tag_reg.tag      = reg2hw.tag_1654.q;
  assign rcache_line[6][118].tag_reg.qe       = reg2hw.tag_1654.qe;
  assign rcache_line[6][118].tag_reg.re       = reg2hw.tag_1654.re;
  assign rcache_line[6][118].status_reg.status = reg2hw.status_1654.q;//status_reg_t'(reg2hw.status_1654.q);
  assign rcache_line[6][118].status_reg.qe    = reg2hw.status_1654.qe;
  assign rcache_line[6][118].status_reg.re    = reg2hw.status_1654.re;


  assign rcache_line[6][119].tag_reg.tag      = reg2hw.tag_1655.q;
  assign rcache_line[6][119].tag_reg.qe       = reg2hw.tag_1655.qe;
  assign rcache_line[6][119].tag_reg.re       = reg2hw.tag_1655.re;
  assign rcache_line[6][119].status_reg.status = reg2hw.status_1655.q;//status_reg_t'(reg2hw.status_1655.q);
  assign rcache_line[6][119].status_reg.qe    = reg2hw.status_1655.qe;
  assign rcache_line[6][119].status_reg.re    = reg2hw.status_1655.re;


  assign rcache_line[6][120].tag_reg.tag      = reg2hw.tag_1656.q;
  assign rcache_line[6][120].tag_reg.qe       = reg2hw.tag_1656.qe;
  assign rcache_line[6][120].tag_reg.re       = reg2hw.tag_1656.re;
  assign rcache_line[6][120].status_reg.status = reg2hw.status_1656.q;//status_reg_t'(reg2hw.status_1656.q);
  assign rcache_line[6][120].status_reg.qe    = reg2hw.status_1656.qe;
  assign rcache_line[6][120].status_reg.re    = reg2hw.status_1656.re;


  assign rcache_line[6][121].tag_reg.tag      = reg2hw.tag_1657.q;
  assign rcache_line[6][121].tag_reg.qe       = reg2hw.tag_1657.qe;
  assign rcache_line[6][121].tag_reg.re       = reg2hw.tag_1657.re;
  assign rcache_line[6][121].status_reg.status = reg2hw.status_1657.q;//status_reg_t'(reg2hw.status_1657.q);
  assign rcache_line[6][121].status_reg.qe    = reg2hw.status_1657.qe;
  assign rcache_line[6][121].status_reg.re    = reg2hw.status_1657.re;


  assign rcache_line[6][122].tag_reg.tag      = reg2hw.tag_1658.q;
  assign rcache_line[6][122].tag_reg.qe       = reg2hw.tag_1658.qe;
  assign rcache_line[6][122].tag_reg.re       = reg2hw.tag_1658.re;
  assign rcache_line[6][122].status_reg.status = reg2hw.status_1658.q;//status_reg_t'(reg2hw.status_1658.q);
  assign rcache_line[6][122].status_reg.qe    = reg2hw.status_1658.qe;
  assign rcache_line[6][122].status_reg.re    = reg2hw.status_1658.re;


  assign rcache_line[6][123].tag_reg.tag      = reg2hw.tag_1659.q;
  assign rcache_line[6][123].tag_reg.qe       = reg2hw.tag_1659.qe;
  assign rcache_line[6][123].tag_reg.re       = reg2hw.tag_1659.re;
  assign rcache_line[6][123].status_reg.status = reg2hw.status_1659.q;//status_reg_t'(reg2hw.status_1659.q);
  assign rcache_line[6][123].status_reg.qe    = reg2hw.status_1659.qe;
  assign rcache_line[6][123].status_reg.re    = reg2hw.status_1659.re;


  assign rcache_line[6][124].tag_reg.tag      = reg2hw.tag_1660.q;
  assign rcache_line[6][124].tag_reg.qe       = reg2hw.tag_1660.qe;
  assign rcache_line[6][124].tag_reg.re       = reg2hw.tag_1660.re;
  assign rcache_line[6][124].status_reg.status = reg2hw.status_1660.q;//status_reg_t'(reg2hw.status_1660.q);
  assign rcache_line[6][124].status_reg.qe    = reg2hw.status_1660.qe;
  assign rcache_line[6][124].status_reg.re    = reg2hw.status_1660.re;


  assign rcache_line[6][125].tag_reg.tag      = reg2hw.tag_1661.q;
  assign rcache_line[6][125].tag_reg.qe       = reg2hw.tag_1661.qe;
  assign rcache_line[6][125].tag_reg.re       = reg2hw.tag_1661.re;
  assign rcache_line[6][125].status_reg.status = reg2hw.status_1661.q;//status_reg_t'(reg2hw.status_1661.q);
  assign rcache_line[6][125].status_reg.qe    = reg2hw.status_1661.qe;
  assign rcache_line[6][125].status_reg.re    = reg2hw.status_1661.re;


  assign rcache_line[6][126].tag_reg.tag      = reg2hw.tag_1662.q;
  assign rcache_line[6][126].tag_reg.qe       = reg2hw.tag_1662.qe;
  assign rcache_line[6][126].tag_reg.re       = reg2hw.tag_1662.re;
  assign rcache_line[6][126].status_reg.status = reg2hw.status_1662.q;//status_reg_t'(reg2hw.status_1662.q);
  assign rcache_line[6][126].status_reg.qe    = reg2hw.status_1662.qe;
  assign rcache_line[6][126].status_reg.re    = reg2hw.status_1662.re;


  assign rcache_line[6][127].tag_reg.tag      = reg2hw.tag_1663.q;
  assign rcache_line[6][127].tag_reg.qe       = reg2hw.tag_1663.qe;
  assign rcache_line[6][127].tag_reg.re       = reg2hw.tag_1663.re;
  assign rcache_line[6][127].status_reg.status = reg2hw.status_1663.q;//status_reg_t'(reg2hw.status_1663.q);
  assign rcache_line[6][127].status_reg.qe    = reg2hw.status_1663.qe;
  assign rcache_line[6][127].status_reg.re    = reg2hw.status_1663.re;


  assign rcache_line[6][128].tag_reg.tag      = reg2hw.tag_1664.q;
  assign rcache_line[6][128].tag_reg.qe       = reg2hw.tag_1664.qe;
  assign rcache_line[6][128].tag_reg.re       = reg2hw.tag_1664.re;
  assign rcache_line[6][128].status_reg.status = reg2hw.status_1664.q;//status_reg_t'(reg2hw.status_1664.q);
  assign rcache_line[6][128].status_reg.qe    = reg2hw.status_1664.qe;
  assign rcache_line[6][128].status_reg.re    = reg2hw.status_1664.re;


  assign rcache_line[6][129].tag_reg.tag      = reg2hw.tag_1665.q;
  assign rcache_line[6][129].tag_reg.qe       = reg2hw.tag_1665.qe;
  assign rcache_line[6][129].tag_reg.re       = reg2hw.tag_1665.re;
  assign rcache_line[6][129].status_reg.status = reg2hw.status_1665.q;//status_reg_t'(reg2hw.status_1665.q);
  assign rcache_line[6][129].status_reg.qe    = reg2hw.status_1665.qe;
  assign rcache_line[6][129].status_reg.re    = reg2hw.status_1665.re;


  assign rcache_line[6][130].tag_reg.tag      = reg2hw.tag_1666.q;
  assign rcache_line[6][130].tag_reg.qe       = reg2hw.tag_1666.qe;
  assign rcache_line[6][130].tag_reg.re       = reg2hw.tag_1666.re;
  assign rcache_line[6][130].status_reg.status = reg2hw.status_1666.q;//status_reg_t'(reg2hw.status_1666.q);
  assign rcache_line[6][130].status_reg.qe    = reg2hw.status_1666.qe;
  assign rcache_line[6][130].status_reg.re    = reg2hw.status_1666.re;


  assign rcache_line[6][131].tag_reg.tag      = reg2hw.tag_1667.q;
  assign rcache_line[6][131].tag_reg.qe       = reg2hw.tag_1667.qe;
  assign rcache_line[6][131].tag_reg.re       = reg2hw.tag_1667.re;
  assign rcache_line[6][131].status_reg.status = reg2hw.status_1667.q;//status_reg_t'(reg2hw.status_1667.q);
  assign rcache_line[6][131].status_reg.qe    = reg2hw.status_1667.qe;
  assign rcache_line[6][131].status_reg.re    = reg2hw.status_1667.re;


  assign rcache_line[6][132].tag_reg.tag      = reg2hw.tag_1668.q;
  assign rcache_line[6][132].tag_reg.qe       = reg2hw.tag_1668.qe;
  assign rcache_line[6][132].tag_reg.re       = reg2hw.tag_1668.re;
  assign rcache_line[6][132].status_reg.status = reg2hw.status_1668.q;//status_reg_t'(reg2hw.status_1668.q);
  assign rcache_line[6][132].status_reg.qe    = reg2hw.status_1668.qe;
  assign rcache_line[6][132].status_reg.re    = reg2hw.status_1668.re;


  assign rcache_line[6][133].tag_reg.tag      = reg2hw.tag_1669.q;
  assign rcache_line[6][133].tag_reg.qe       = reg2hw.tag_1669.qe;
  assign rcache_line[6][133].tag_reg.re       = reg2hw.tag_1669.re;
  assign rcache_line[6][133].status_reg.status = reg2hw.status_1669.q;//status_reg_t'(reg2hw.status_1669.q);
  assign rcache_line[6][133].status_reg.qe    = reg2hw.status_1669.qe;
  assign rcache_line[6][133].status_reg.re    = reg2hw.status_1669.re;


  assign rcache_line[6][134].tag_reg.tag      = reg2hw.tag_1670.q;
  assign rcache_line[6][134].tag_reg.qe       = reg2hw.tag_1670.qe;
  assign rcache_line[6][134].tag_reg.re       = reg2hw.tag_1670.re;
  assign rcache_line[6][134].status_reg.status = reg2hw.status_1670.q;//status_reg_t'(reg2hw.status_1670.q);
  assign rcache_line[6][134].status_reg.qe    = reg2hw.status_1670.qe;
  assign rcache_line[6][134].status_reg.re    = reg2hw.status_1670.re;


  assign rcache_line[6][135].tag_reg.tag      = reg2hw.tag_1671.q;
  assign rcache_line[6][135].tag_reg.qe       = reg2hw.tag_1671.qe;
  assign rcache_line[6][135].tag_reg.re       = reg2hw.tag_1671.re;
  assign rcache_line[6][135].status_reg.status = reg2hw.status_1671.q;//status_reg_t'(reg2hw.status_1671.q);
  assign rcache_line[6][135].status_reg.qe    = reg2hw.status_1671.qe;
  assign rcache_line[6][135].status_reg.re    = reg2hw.status_1671.re;


  assign rcache_line[6][136].tag_reg.tag      = reg2hw.tag_1672.q;
  assign rcache_line[6][136].tag_reg.qe       = reg2hw.tag_1672.qe;
  assign rcache_line[6][136].tag_reg.re       = reg2hw.tag_1672.re;
  assign rcache_line[6][136].status_reg.status = reg2hw.status_1672.q;//status_reg_t'(reg2hw.status_1672.q);
  assign rcache_line[6][136].status_reg.qe    = reg2hw.status_1672.qe;
  assign rcache_line[6][136].status_reg.re    = reg2hw.status_1672.re;


  assign rcache_line[6][137].tag_reg.tag      = reg2hw.tag_1673.q;
  assign rcache_line[6][137].tag_reg.qe       = reg2hw.tag_1673.qe;
  assign rcache_line[6][137].tag_reg.re       = reg2hw.tag_1673.re;
  assign rcache_line[6][137].status_reg.status = reg2hw.status_1673.q;//status_reg_t'(reg2hw.status_1673.q);
  assign rcache_line[6][137].status_reg.qe    = reg2hw.status_1673.qe;
  assign rcache_line[6][137].status_reg.re    = reg2hw.status_1673.re;


  assign rcache_line[6][138].tag_reg.tag      = reg2hw.tag_1674.q;
  assign rcache_line[6][138].tag_reg.qe       = reg2hw.tag_1674.qe;
  assign rcache_line[6][138].tag_reg.re       = reg2hw.tag_1674.re;
  assign rcache_line[6][138].status_reg.status = reg2hw.status_1674.q;//status_reg_t'(reg2hw.status_1674.q);
  assign rcache_line[6][138].status_reg.qe    = reg2hw.status_1674.qe;
  assign rcache_line[6][138].status_reg.re    = reg2hw.status_1674.re;


  assign rcache_line[6][139].tag_reg.tag      = reg2hw.tag_1675.q;
  assign rcache_line[6][139].tag_reg.qe       = reg2hw.tag_1675.qe;
  assign rcache_line[6][139].tag_reg.re       = reg2hw.tag_1675.re;
  assign rcache_line[6][139].status_reg.status = reg2hw.status_1675.q;//status_reg_t'(reg2hw.status_1675.q);
  assign rcache_line[6][139].status_reg.qe    = reg2hw.status_1675.qe;
  assign rcache_line[6][139].status_reg.re    = reg2hw.status_1675.re;


  assign rcache_line[6][140].tag_reg.tag      = reg2hw.tag_1676.q;
  assign rcache_line[6][140].tag_reg.qe       = reg2hw.tag_1676.qe;
  assign rcache_line[6][140].tag_reg.re       = reg2hw.tag_1676.re;
  assign rcache_line[6][140].status_reg.status = reg2hw.status_1676.q;//status_reg_t'(reg2hw.status_1676.q);
  assign rcache_line[6][140].status_reg.qe    = reg2hw.status_1676.qe;
  assign rcache_line[6][140].status_reg.re    = reg2hw.status_1676.re;


  assign rcache_line[6][141].tag_reg.tag      = reg2hw.tag_1677.q;
  assign rcache_line[6][141].tag_reg.qe       = reg2hw.tag_1677.qe;
  assign rcache_line[6][141].tag_reg.re       = reg2hw.tag_1677.re;
  assign rcache_line[6][141].status_reg.status = reg2hw.status_1677.q;//status_reg_t'(reg2hw.status_1677.q);
  assign rcache_line[6][141].status_reg.qe    = reg2hw.status_1677.qe;
  assign rcache_line[6][141].status_reg.re    = reg2hw.status_1677.re;


  assign rcache_line[6][142].tag_reg.tag      = reg2hw.tag_1678.q;
  assign rcache_line[6][142].tag_reg.qe       = reg2hw.tag_1678.qe;
  assign rcache_line[6][142].tag_reg.re       = reg2hw.tag_1678.re;
  assign rcache_line[6][142].status_reg.status = reg2hw.status_1678.q;//status_reg_t'(reg2hw.status_1678.q);
  assign rcache_line[6][142].status_reg.qe    = reg2hw.status_1678.qe;
  assign rcache_line[6][142].status_reg.re    = reg2hw.status_1678.re;


  assign rcache_line[6][143].tag_reg.tag      = reg2hw.tag_1679.q;
  assign rcache_line[6][143].tag_reg.qe       = reg2hw.tag_1679.qe;
  assign rcache_line[6][143].tag_reg.re       = reg2hw.tag_1679.re;
  assign rcache_line[6][143].status_reg.status = reg2hw.status_1679.q;//status_reg_t'(reg2hw.status_1679.q);
  assign rcache_line[6][143].status_reg.qe    = reg2hw.status_1679.qe;
  assign rcache_line[6][143].status_reg.re    = reg2hw.status_1679.re;


  assign rcache_line[6][144].tag_reg.tag      = reg2hw.tag_1680.q;
  assign rcache_line[6][144].tag_reg.qe       = reg2hw.tag_1680.qe;
  assign rcache_line[6][144].tag_reg.re       = reg2hw.tag_1680.re;
  assign rcache_line[6][144].status_reg.status = reg2hw.status_1680.q;//status_reg_t'(reg2hw.status_1680.q);
  assign rcache_line[6][144].status_reg.qe    = reg2hw.status_1680.qe;
  assign rcache_line[6][144].status_reg.re    = reg2hw.status_1680.re;


  assign rcache_line[6][145].tag_reg.tag      = reg2hw.tag_1681.q;
  assign rcache_line[6][145].tag_reg.qe       = reg2hw.tag_1681.qe;
  assign rcache_line[6][145].tag_reg.re       = reg2hw.tag_1681.re;
  assign rcache_line[6][145].status_reg.status = reg2hw.status_1681.q;//status_reg_t'(reg2hw.status_1681.q);
  assign rcache_line[6][145].status_reg.qe    = reg2hw.status_1681.qe;
  assign rcache_line[6][145].status_reg.re    = reg2hw.status_1681.re;


  assign rcache_line[6][146].tag_reg.tag      = reg2hw.tag_1682.q;
  assign rcache_line[6][146].tag_reg.qe       = reg2hw.tag_1682.qe;
  assign rcache_line[6][146].tag_reg.re       = reg2hw.tag_1682.re;
  assign rcache_line[6][146].status_reg.status = reg2hw.status_1682.q;//status_reg_t'(reg2hw.status_1682.q);
  assign rcache_line[6][146].status_reg.qe    = reg2hw.status_1682.qe;
  assign rcache_line[6][146].status_reg.re    = reg2hw.status_1682.re;


  assign rcache_line[6][147].tag_reg.tag      = reg2hw.tag_1683.q;
  assign rcache_line[6][147].tag_reg.qe       = reg2hw.tag_1683.qe;
  assign rcache_line[6][147].tag_reg.re       = reg2hw.tag_1683.re;
  assign rcache_line[6][147].status_reg.status = reg2hw.status_1683.q;//status_reg_t'(reg2hw.status_1683.q);
  assign rcache_line[6][147].status_reg.qe    = reg2hw.status_1683.qe;
  assign rcache_line[6][147].status_reg.re    = reg2hw.status_1683.re;


  assign rcache_line[6][148].tag_reg.tag      = reg2hw.tag_1684.q;
  assign rcache_line[6][148].tag_reg.qe       = reg2hw.tag_1684.qe;
  assign rcache_line[6][148].tag_reg.re       = reg2hw.tag_1684.re;
  assign rcache_line[6][148].status_reg.status = reg2hw.status_1684.q;//status_reg_t'(reg2hw.status_1684.q);
  assign rcache_line[6][148].status_reg.qe    = reg2hw.status_1684.qe;
  assign rcache_line[6][148].status_reg.re    = reg2hw.status_1684.re;


  assign rcache_line[6][149].tag_reg.tag      = reg2hw.tag_1685.q;
  assign rcache_line[6][149].tag_reg.qe       = reg2hw.tag_1685.qe;
  assign rcache_line[6][149].tag_reg.re       = reg2hw.tag_1685.re;
  assign rcache_line[6][149].status_reg.status = reg2hw.status_1685.q;//status_reg_t'(reg2hw.status_1685.q);
  assign rcache_line[6][149].status_reg.qe    = reg2hw.status_1685.qe;
  assign rcache_line[6][149].status_reg.re    = reg2hw.status_1685.re;


  assign rcache_line[6][150].tag_reg.tag      = reg2hw.tag_1686.q;
  assign rcache_line[6][150].tag_reg.qe       = reg2hw.tag_1686.qe;
  assign rcache_line[6][150].tag_reg.re       = reg2hw.tag_1686.re;
  assign rcache_line[6][150].status_reg.status = reg2hw.status_1686.q;//status_reg_t'(reg2hw.status_1686.q);
  assign rcache_line[6][150].status_reg.qe    = reg2hw.status_1686.qe;
  assign rcache_line[6][150].status_reg.re    = reg2hw.status_1686.re;


  assign rcache_line[6][151].tag_reg.tag      = reg2hw.tag_1687.q;
  assign rcache_line[6][151].tag_reg.qe       = reg2hw.tag_1687.qe;
  assign rcache_line[6][151].tag_reg.re       = reg2hw.tag_1687.re;
  assign rcache_line[6][151].status_reg.status = reg2hw.status_1687.q;//status_reg_t'(reg2hw.status_1687.q);
  assign rcache_line[6][151].status_reg.qe    = reg2hw.status_1687.qe;
  assign rcache_line[6][151].status_reg.re    = reg2hw.status_1687.re;


  assign rcache_line[6][152].tag_reg.tag      = reg2hw.tag_1688.q;
  assign rcache_line[6][152].tag_reg.qe       = reg2hw.tag_1688.qe;
  assign rcache_line[6][152].tag_reg.re       = reg2hw.tag_1688.re;
  assign rcache_line[6][152].status_reg.status = reg2hw.status_1688.q;//status_reg_t'(reg2hw.status_1688.q);
  assign rcache_line[6][152].status_reg.qe    = reg2hw.status_1688.qe;
  assign rcache_line[6][152].status_reg.re    = reg2hw.status_1688.re;


  assign rcache_line[6][153].tag_reg.tag      = reg2hw.tag_1689.q;
  assign rcache_line[6][153].tag_reg.qe       = reg2hw.tag_1689.qe;
  assign rcache_line[6][153].tag_reg.re       = reg2hw.tag_1689.re;
  assign rcache_line[6][153].status_reg.status = reg2hw.status_1689.q;//status_reg_t'(reg2hw.status_1689.q);
  assign rcache_line[6][153].status_reg.qe    = reg2hw.status_1689.qe;
  assign rcache_line[6][153].status_reg.re    = reg2hw.status_1689.re;


  assign rcache_line[6][154].tag_reg.tag      = reg2hw.tag_1690.q;
  assign rcache_line[6][154].tag_reg.qe       = reg2hw.tag_1690.qe;
  assign rcache_line[6][154].tag_reg.re       = reg2hw.tag_1690.re;
  assign rcache_line[6][154].status_reg.status = reg2hw.status_1690.q;//status_reg_t'(reg2hw.status_1690.q);
  assign rcache_line[6][154].status_reg.qe    = reg2hw.status_1690.qe;
  assign rcache_line[6][154].status_reg.re    = reg2hw.status_1690.re;


  assign rcache_line[6][155].tag_reg.tag      = reg2hw.tag_1691.q;
  assign rcache_line[6][155].tag_reg.qe       = reg2hw.tag_1691.qe;
  assign rcache_line[6][155].tag_reg.re       = reg2hw.tag_1691.re;
  assign rcache_line[6][155].status_reg.status = reg2hw.status_1691.q;//status_reg_t'(reg2hw.status_1691.q);
  assign rcache_line[6][155].status_reg.qe    = reg2hw.status_1691.qe;
  assign rcache_line[6][155].status_reg.re    = reg2hw.status_1691.re;


  assign rcache_line[6][156].tag_reg.tag      = reg2hw.tag_1692.q;
  assign rcache_line[6][156].tag_reg.qe       = reg2hw.tag_1692.qe;
  assign rcache_line[6][156].tag_reg.re       = reg2hw.tag_1692.re;
  assign rcache_line[6][156].status_reg.status = reg2hw.status_1692.q;//status_reg_t'(reg2hw.status_1692.q);
  assign rcache_line[6][156].status_reg.qe    = reg2hw.status_1692.qe;
  assign rcache_line[6][156].status_reg.re    = reg2hw.status_1692.re;


  assign rcache_line[6][157].tag_reg.tag      = reg2hw.tag_1693.q;
  assign rcache_line[6][157].tag_reg.qe       = reg2hw.tag_1693.qe;
  assign rcache_line[6][157].tag_reg.re       = reg2hw.tag_1693.re;
  assign rcache_line[6][157].status_reg.status = reg2hw.status_1693.q;//status_reg_t'(reg2hw.status_1693.q);
  assign rcache_line[6][157].status_reg.qe    = reg2hw.status_1693.qe;
  assign rcache_line[6][157].status_reg.re    = reg2hw.status_1693.re;


  assign rcache_line[6][158].tag_reg.tag      = reg2hw.tag_1694.q;
  assign rcache_line[6][158].tag_reg.qe       = reg2hw.tag_1694.qe;
  assign rcache_line[6][158].tag_reg.re       = reg2hw.tag_1694.re;
  assign rcache_line[6][158].status_reg.status = reg2hw.status_1694.q;//status_reg_t'(reg2hw.status_1694.q);
  assign rcache_line[6][158].status_reg.qe    = reg2hw.status_1694.qe;
  assign rcache_line[6][158].status_reg.re    = reg2hw.status_1694.re;


  assign rcache_line[6][159].tag_reg.tag      = reg2hw.tag_1695.q;
  assign rcache_line[6][159].tag_reg.qe       = reg2hw.tag_1695.qe;
  assign rcache_line[6][159].tag_reg.re       = reg2hw.tag_1695.re;
  assign rcache_line[6][159].status_reg.status = reg2hw.status_1695.q;//status_reg_t'(reg2hw.status_1695.q);
  assign rcache_line[6][159].status_reg.qe    = reg2hw.status_1695.qe;
  assign rcache_line[6][159].status_reg.re    = reg2hw.status_1695.re;


  assign rcache_line[6][160].tag_reg.tag      = reg2hw.tag_1696.q;
  assign rcache_line[6][160].tag_reg.qe       = reg2hw.tag_1696.qe;
  assign rcache_line[6][160].tag_reg.re       = reg2hw.tag_1696.re;
  assign rcache_line[6][160].status_reg.status = reg2hw.status_1696.q;//status_reg_t'(reg2hw.status_1696.q);
  assign rcache_line[6][160].status_reg.qe    = reg2hw.status_1696.qe;
  assign rcache_line[6][160].status_reg.re    = reg2hw.status_1696.re;


  assign rcache_line[6][161].tag_reg.tag      = reg2hw.tag_1697.q;
  assign rcache_line[6][161].tag_reg.qe       = reg2hw.tag_1697.qe;
  assign rcache_line[6][161].tag_reg.re       = reg2hw.tag_1697.re;
  assign rcache_line[6][161].status_reg.status = reg2hw.status_1697.q;//status_reg_t'(reg2hw.status_1697.q);
  assign rcache_line[6][161].status_reg.qe    = reg2hw.status_1697.qe;
  assign rcache_line[6][161].status_reg.re    = reg2hw.status_1697.re;


  assign rcache_line[6][162].tag_reg.tag      = reg2hw.tag_1698.q;
  assign rcache_line[6][162].tag_reg.qe       = reg2hw.tag_1698.qe;
  assign rcache_line[6][162].tag_reg.re       = reg2hw.tag_1698.re;
  assign rcache_line[6][162].status_reg.status = reg2hw.status_1698.q;//status_reg_t'(reg2hw.status_1698.q);
  assign rcache_line[6][162].status_reg.qe    = reg2hw.status_1698.qe;
  assign rcache_line[6][162].status_reg.re    = reg2hw.status_1698.re;


  assign rcache_line[6][163].tag_reg.tag      = reg2hw.tag_1699.q;
  assign rcache_line[6][163].tag_reg.qe       = reg2hw.tag_1699.qe;
  assign rcache_line[6][163].tag_reg.re       = reg2hw.tag_1699.re;
  assign rcache_line[6][163].status_reg.status = reg2hw.status_1699.q;//status_reg_t'(reg2hw.status_1699.q);
  assign rcache_line[6][163].status_reg.qe    = reg2hw.status_1699.qe;
  assign rcache_line[6][163].status_reg.re    = reg2hw.status_1699.re;


  assign rcache_line[6][164].tag_reg.tag      = reg2hw.tag_1700.q;
  assign rcache_line[6][164].tag_reg.qe       = reg2hw.tag_1700.qe;
  assign rcache_line[6][164].tag_reg.re       = reg2hw.tag_1700.re;
  assign rcache_line[6][164].status_reg.status = reg2hw.status_1700.q;//status_reg_t'(reg2hw.status_1700.q);
  assign rcache_line[6][164].status_reg.qe    = reg2hw.status_1700.qe;
  assign rcache_line[6][164].status_reg.re    = reg2hw.status_1700.re;


  assign rcache_line[6][165].tag_reg.tag      = reg2hw.tag_1701.q;
  assign rcache_line[6][165].tag_reg.qe       = reg2hw.tag_1701.qe;
  assign rcache_line[6][165].tag_reg.re       = reg2hw.tag_1701.re;
  assign rcache_line[6][165].status_reg.status = reg2hw.status_1701.q;//status_reg_t'(reg2hw.status_1701.q);
  assign rcache_line[6][165].status_reg.qe    = reg2hw.status_1701.qe;
  assign rcache_line[6][165].status_reg.re    = reg2hw.status_1701.re;


  assign rcache_line[6][166].tag_reg.tag      = reg2hw.tag_1702.q;
  assign rcache_line[6][166].tag_reg.qe       = reg2hw.tag_1702.qe;
  assign rcache_line[6][166].tag_reg.re       = reg2hw.tag_1702.re;
  assign rcache_line[6][166].status_reg.status = reg2hw.status_1702.q;//status_reg_t'(reg2hw.status_1702.q);
  assign rcache_line[6][166].status_reg.qe    = reg2hw.status_1702.qe;
  assign rcache_line[6][166].status_reg.re    = reg2hw.status_1702.re;


  assign rcache_line[6][167].tag_reg.tag      = reg2hw.tag_1703.q;
  assign rcache_line[6][167].tag_reg.qe       = reg2hw.tag_1703.qe;
  assign rcache_line[6][167].tag_reg.re       = reg2hw.tag_1703.re;
  assign rcache_line[6][167].status_reg.status = reg2hw.status_1703.q;//status_reg_t'(reg2hw.status_1703.q);
  assign rcache_line[6][167].status_reg.qe    = reg2hw.status_1703.qe;
  assign rcache_line[6][167].status_reg.re    = reg2hw.status_1703.re;


  assign rcache_line[6][168].tag_reg.tag      = reg2hw.tag_1704.q;
  assign rcache_line[6][168].tag_reg.qe       = reg2hw.tag_1704.qe;
  assign rcache_line[6][168].tag_reg.re       = reg2hw.tag_1704.re;
  assign rcache_line[6][168].status_reg.status = reg2hw.status_1704.q;//status_reg_t'(reg2hw.status_1704.q);
  assign rcache_line[6][168].status_reg.qe    = reg2hw.status_1704.qe;
  assign rcache_line[6][168].status_reg.re    = reg2hw.status_1704.re;


  assign rcache_line[6][169].tag_reg.tag      = reg2hw.tag_1705.q;
  assign rcache_line[6][169].tag_reg.qe       = reg2hw.tag_1705.qe;
  assign rcache_line[6][169].tag_reg.re       = reg2hw.tag_1705.re;
  assign rcache_line[6][169].status_reg.status = reg2hw.status_1705.q;//status_reg_t'(reg2hw.status_1705.q);
  assign rcache_line[6][169].status_reg.qe    = reg2hw.status_1705.qe;
  assign rcache_line[6][169].status_reg.re    = reg2hw.status_1705.re;


  assign rcache_line[6][170].tag_reg.tag      = reg2hw.tag_1706.q;
  assign rcache_line[6][170].tag_reg.qe       = reg2hw.tag_1706.qe;
  assign rcache_line[6][170].tag_reg.re       = reg2hw.tag_1706.re;
  assign rcache_line[6][170].status_reg.status = reg2hw.status_1706.q;//status_reg_t'(reg2hw.status_1706.q);
  assign rcache_line[6][170].status_reg.qe    = reg2hw.status_1706.qe;
  assign rcache_line[6][170].status_reg.re    = reg2hw.status_1706.re;


  assign rcache_line[6][171].tag_reg.tag      = reg2hw.tag_1707.q;
  assign rcache_line[6][171].tag_reg.qe       = reg2hw.tag_1707.qe;
  assign rcache_line[6][171].tag_reg.re       = reg2hw.tag_1707.re;
  assign rcache_line[6][171].status_reg.status = reg2hw.status_1707.q;//status_reg_t'(reg2hw.status_1707.q);
  assign rcache_line[6][171].status_reg.qe    = reg2hw.status_1707.qe;
  assign rcache_line[6][171].status_reg.re    = reg2hw.status_1707.re;


  assign rcache_line[6][172].tag_reg.tag      = reg2hw.tag_1708.q;
  assign rcache_line[6][172].tag_reg.qe       = reg2hw.tag_1708.qe;
  assign rcache_line[6][172].tag_reg.re       = reg2hw.tag_1708.re;
  assign rcache_line[6][172].status_reg.status = reg2hw.status_1708.q;//status_reg_t'(reg2hw.status_1708.q);
  assign rcache_line[6][172].status_reg.qe    = reg2hw.status_1708.qe;
  assign rcache_line[6][172].status_reg.re    = reg2hw.status_1708.re;


  assign rcache_line[6][173].tag_reg.tag      = reg2hw.tag_1709.q;
  assign rcache_line[6][173].tag_reg.qe       = reg2hw.tag_1709.qe;
  assign rcache_line[6][173].tag_reg.re       = reg2hw.tag_1709.re;
  assign rcache_line[6][173].status_reg.status = reg2hw.status_1709.q;//status_reg_t'(reg2hw.status_1709.q);
  assign rcache_line[6][173].status_reg.qe    = reg2hw.status_1709.qe;
  assign rcache_line[6][173].status_reg.re    = reg2hw.status_1709.re;


  assign rcache_line[6][174].tag_reg.tag      = reg2hw.tag_1710.q;
  assign rcache_line[6][174].tag_reg.qe       = reg2hw.tag_1710.qe;
  assign rcache_line[6][174].tag_reg.re       = reg2hw.tag_1710.re;
  assign rcache_line[6][174].status_reg.status = reg2hw.status_1710.q;//status_reg_t'(reg2hw.status_1710.q);
  assign rcache_line[6][174].status_reg.qe    = reg2hw.status_1710.qe;
  assign rcache_line[6][174].status_reg.re    = reg2hw.status_1710.re;


  assign rcache_line[6][175].tag_reg.tag      = reg2hw.tag_1711.q;
  assign rcache_line[6][175].tag_reg.qe       = reg2hw.tag_1711.qe;
  assign rcache_line[6][175].tag_reg.re       = reg2hw.tag_1711.re;
  assign rcache_line[6][175].status_reg.status = reg2hw.status_1711.q;//status_reg_t'(reg2hw.status_1711.q);
  assign rcache_line[6][175].status_reg.qe    = reg2hw.status_1711.qe;
  assign rcache_line[6][175].status_reg.re    = reg2hw.status_1711.re;


  assign rcache_line[6][176].tag_reg.tag      = reg2hw.tag_1712.q;
  assign rcache_line[6][176].tag_reg.qe       = reg2hw.tag_1712.qe;
  assign rcache_line[6][176].tag_reg.re       = reg2hw.tag_1712.re;
  assign rcache_line[6][176].status_reg.status = reg2hw.status_1712.q;//status_reg_t'(reg2hw.status_1712.q);
  assign rcache_line[6][176].status_reg.qe    = reg2hw.status_1712.qe;
  assign rcache_line[6][176].status_reg.re    = reg2hw.status_1712.re;


  assign rcache_line[6][177].tag_reg.tag      = reg2hw.tag_1713.q;
  assign rcache_line[6][177].tag_reg.qe       = reg2hw.tag_1713.qe;
  assign rcache_line[6][177].tag_reg.re       = reg2hw.tag_1713.re;
  assign rcache_line[6][177].status_reg.status = reg2hw.status_1713.q;//status_reg_t'(reg2hw.status_1713.q);
  assign rcache_line[6][177].status_reg.qe    = reg2hw.status_1713.qe;
  assign rcache_line[6][177].status_reg.re    = reg2hw.status_1713.re;


  assign rcache_line[6][178].tag_reg.tag      = reg2hw.tag_1714.q;
  assign rcache_line[6][178].tag_reg.qe       = reg2hw.tag_1714.qe;
  assign rcache_line[6][178].tag_reg.re       = reg2hw.tag_1714.re;
  assign rcache_line[6][178].status_reg.status = reg2hw.status_1714.q;//status_reg_t'(reg2hw.status_1714.q);
  assign rcache_line[6][178].status_reg.qe    = reg2hw.status_1714.qe;
  assign rcache_line[6][178].status_reg.re    = reg2hw.status_1714.re;


  assign rcache_line[6][179].tag_reg.tag      = reg2hw.tag_1715.q;
  assign rcache_line[6][179].tag_reg.qe       = reg2hw.tag_1715.qe;
  assign rcache_line[6][179].tag_reg.re       = reg2hw.tag_1715.re;
  assign rcache_line[6][179].status_reg.status = reg2hw.status_1715.q;//status_reg_t'(reg2hw.status_1715.q);
  assign rcache_line[6][179].status_reg.qe    = reg2hw.status_1715.qe;
  assign rcache_line[6][179].status_reg.re    = reg2hw.status_1715.re;


  assign rcache_line[6][180].tag_reg.tag      = reg2hw.tag_1716.q;
  assign rcache_line[6][180].tag_reg.qe       = reg2hw.tag_1716.qe;
  assign rcache_line[6][180].tag_reg.re       = reg2hw.tag_1716.re;
  assign rcache_line[6][180].status_reg.status = reg2hw.status_1716.q;//status_reg_t'(reg2hw.status_1716.q);
  assign rcache_line[6][180].status_reg.qe    = reg2hw.status_1716.qe;
  assign rcache_line[6][180].status_reg.re    = reg2hw.status_1716.re;


  assign rcache_line[6][181].tag_reg.tag      = reg2hw.tag_1717.q;
  assign rcache_line[6][181].tag_reg.qe       = reg2hw.tag_1717.qe;
  assign rcache_line[6][181].tag_reg.re       = reg2hw.tag_1717.re;
  assign rcache_line[6][181].status_reg.status = reg2hw.status_1717.q;//status_reg_t'(reg2hw.status_1717.q);
  assign rcache_line[6][181].status_reg.qe    = reg2hw.status_1717.qe;
  assign rcache_line[6][181].status_reg.re    = reg2hw.status_1717.re;


  assign rcache_line[6][182].tag_reg.tag      = reg2hw.tag_1718.q;
  assign rcache_line[6][182].tag_reg.qe       = reg2hw.tag_1718.qe;
  assign rcache_line[6][182].tag_reg.re       = reg2hw.tag_1718.re;
  assign rcache_line[6][182].status_reg.status = reg2hw.status_1718.q;//status_reg_t'(reg2hw.status_1718.q);
  assign rcache_line[6][182].status_reg.qe    = reg2hw.status_1718.qe;
  assign rcache_line[6][182].status_reg.re    = reg2hw.status_1718.re;


  assign rcache_line[6][183].tag_reg.tag      = reg2hw.tag_1719.q;
  assign rcache_line[6][183].tag_reg.qe       = reg2hw.tag_1719.qe;
  assign rcache_line[6][183].tag_reg.re       = reg2hw.tag_1719.re;
  assign rcache_line[6][183].status_reg.status = reg2hw.status_1719.q;//status_reg_t'(reg2hw.status_1719.q);
  assign rcache_line[6][183].status_reg.qe    = reg2hw.status_1719.qe;
  assign rcache_line[6][183].status_reg.re    = reg2hw.status_1719.re;


  assign rcache_line[6][184].tag_reg.tag      = reg2hw.tag_1720.q;
  assign rcache_line[6][184].tag_reg.qe       = reg2hw.tag_1720.qe;
  assign rcache_line[6][184].tag_reg.re       = reg2hw.tag_1720.re;
  assign rcache_line[6][184].status_reg.status = reg2hw.status_1720.q;//status_reg_t'(reg2hw.status_1720.q);
  assign rcache_line[6][184].status_reg.qe    = reg2hw.status_1720.qe;
  assign rcache_line[6][184].status_reg.re    = reg2hw.status_1720.re;


  assign rcache_line[6][185].tag_reg.tag      = reg2hw.tag_1721.q;
  assign rcache_line[6][185].tag_reg.qe       = reg2hw.tag_1721.qe;
  assign rcache_line[6][185].tag_reg.re       = reg2hw.tag_1721.re;
  assign rcache_line[6][185].status_reg.status = reg2hw.status_1721.q;//status_reg_t'(reg2hw.status_1721.q);
  assign rcache_line[6][185].status_reg.qe    = reg2hw.status_1721.qe;
  assign rcache_line[6][185].status_reg.re    = reg2hw.status_1721.re;


  assign rcache_line[6][186].tag_reg.tag      = reg2hw.tag_1722.q;
  assign rcache_line[6][186].tag_reg.qe       = reg2hw.tag_1722.qe;
  assign rcache_line[6][186].tag_reg.re       = reg2hw.tag_1722.re;
  assign rcache_line[6][186].status_reg.status = reg2hw.status_1722.q;//status_reg_t'(reg2hw.status_1722.q);
  assign rcache_line[6][186].status_reg.qe    = reg2hw.status_1722.qe;
  assign rcache_line[6][186].status_reg.re    = reg2hw.status_1722.re;


  assign rcache_line[6][187].tag_reg.tag      = reg2hw.tag_1723.q;
  assign rcache_line[6][187].tag_reg.qe       = reg2hw.tag_1723.qe;
  assign rcache_line[6][187].tag_reg.re       = reg2hw.tag_1723.re;
  assign rcache_line[6][187].status_reg.status = reg2hw.status_1723.q;//status_reg_t'(reg2hw.status_1723.q);
  assign rcache_line[6][187].status_reg.qe    = reg2hw.status_1723.qe;
  assign rcache_line[6][187].status_reg.re    = reg2hw.status_1723.re;


  assign rcache_line[6][188].tag_reg.tag      = reg2hw.tag_1724.q;
  assign rcache_line[6][188].tag_reg.qe       = reg2hw.tag_1724.qe;
  assign rcache_line[6][188].tag_reg.re       = reg2hw.tag_1724.re;
  assign rcache_line[6][188].status_reg.status = reg2hw.status_1724.q;//status_reg_t'(reg2hw.status_1724.q);
  assign rcache_line[6][188].status_reg.qe    = reg2hw.status_1724.qe;
  assign rcache_line[6][188].status_reg.re    = reg2hw.status_1724.re;


  assign rcache_line[6][189].tag_reg.tag      = reg2hw.tag_1725.q;
  assign rcache_line[6][189].tag_reg.qe       = reg2hw.tag_1725.qe;
  assign rcache_line[6][189].tag_reg.re       = reg2hw.tag_1725.re;
  assign rcache_line[6][189].status_reg.status = reg2hw.status_1725.q;//status_reg_t'(reg2hw.status_1725.q);
  assign rcache_line[6][189].status_reg.qe    = reg2hw.status_1725.qe;
  assign rcache_line[6][189].status_reg.re    = reg2hw.status_1725.re;


  assign rcache_line[6][190].tag_reg.tag      = reg2hw.tag_1726.q;
  assign rcache_line[6][190].tag_reg.qe       = reg2hw.tag_1726.qe;
  assign rcache_line[6][190].tag_reg.re       = reg2hw.tag_1726.re;
  assign rcache_line[6][190].status_reg.status = reg2hw.status_1726.q;//status_reg_t'(reg2hw.status_1726.q);
  assign rcache_line[6][190].status_reg.qe    = reg2hw.status_1726.qe;
  assign rcache_line[6][190].status_reg.re    = reg2hw.status_1726.re;


  assign rcache_line[6][191].tag_reg.tag      = reg2hw.tag_1727.q;
  assign rcache_line[6][191].tag_reg.qe       = reg2hw.tag_1727.qe;
  assign rcache_line[6][191].tag_reg.re       = reg2hw.tag_1727.re;
  assign rcache_line[6][191].status_reg.status = reg2hw.status_1727.q;//status_reg_t'(reg2hw.status_1727.q);
  assign rcache_line[6][191].status_reg.qe    = reg2hw.status_1727.qe;
  assign rcache_line[6][191].status_reg.re    = reg2hw.status_1727.re;


  assign rcache_line[6][192].tag_reg.tag      = reg2hw.tag_1728.q;
  assign rcache_line[6][192].tag_reg.qe       = reg2hw.tag_1728.qe;
  assign rcache_line[6][192].tag_reg.re       = reg2hw.tag_1728.re;
  assign rcache_line[6][192].status_reg.status = reg2hw.status_1728.q;//status_reg_t'(reg2hw.status_1728.q);
  assign rcache_line[6][192].status_reg.qe    = reg2hw.status_1728.qe;
  assign rcache_line[6][192].status_reg.re    = reg2hw.status_1728.re;


  assign rcache_line[6][193].tag_reg.tag      = reg2hw.tag_1729.q;
  assign rcache_line[6][193].tag_reg.qe       = reg2hw.tag_1729.qe;
  assign rcache_line[6][193].tag_reg.re       = reg2hw.tag_1729.re;
  assign rcache_line[6][193].status_reg.status = reg2hw.status_1729.q;//status_reg_t'(reg2hw.status_1729.q);
  assign rcache_line[6][193].status_reg.qe    = reg2hw.status_1729.qe;
  assign rcache_line[6][193].status_reg.re    = reg2hw.status_1729.re;


  assign rcache_line[6][194].tag_reg.tag      = reg2hw.tag_1730.q;
  assign rcache_line[6][194].tag_reg.qe       = reg2hw.tag_1730.qe;
  assign rcache_line[6][194].tag_reg.re       = reg2hw.tag_1730.re;
  assign rcache_line[6][194].status_reg.status = reg2hw.status_1730.q;//status_reg_t'(reg2hw.status_1730.q);
  assign rcache_line[6][194].status_reg.qe    = reg2hw.status_1730.qe;
  assign rcache_line[6][194].status_reg.re    = reg2hw.status_1730.re;


  assign rcache_line[6][195].tag_reg.tag      = reg2hw.tag_1731.q;
  assign rcache_line[6][195].tag_reg.qe       = reg2hw.tag_1731.qe;
  assign rcache_line[6][195].tag_reg.re       = reg2hw.tag_1731.re;
  assign rcache_line[6][195].status_reg.status = reg2hw.status_1731.q;//status_reg_t'(reg2hw.status_1731.q);
  assign rcache_line[6][195].status_reg.qe    = reg2hw.status_1731.qe;
  assign rcache_line[6][195].status_reg.re    = reg2hw.status_1731.re;


  assign rcache_line[6][196].tag_reg.tag      = reg2hw.tag_1732.q;
  assign rcache_line[6][196].tag_reg.qe       = reg2hw.tag_1732.qe;
  assign rcache_line[6][196].tag_reg.re       = reg2hw.tag_1732.re;
  assign rcache_line[6][196].status_reg.status = reg2hw.status_1732.q;//status_reg_t'(reg2hw.status_1732.q);
  assign rcache_line[6][196].status_reg.qe    = reg2hw.status_1732.qe;
  assign rcache_line[6][196].status_reg.re    = reg2hw.status_1732.re;


  assign rcache_line[6][197].tag_reg.tag      = reg2hw.tag_1733.q;
  assign rcache_line[6][197].tag_reg.qe       = reg2hw.tag_1733.qe;
  assign rcache_line[6][197].tag_reg.re       = reg2hw.tag_1733.re;
  assign rcache_line[6][197].status_reg.status = reg2hw.status_1733.q;//status_reg_t'(reg2hw.status_1733.q);
  assign rcache_line[6][197].status_reg.qe    = reg2hw.status_1733.qe;
  assign rcache_line[6][197].status_reg.re    = reg2hw.status_1733.re;


  assign rcache_line[6][198].tag_reg.tag      = reg2hw.tag_1734.q;
  assign rcache_line[6][198].tag_reg.qe       = reg2hw.tag_1734.qe;
  assign rcache_line[6][198].tag_reg.re       = reg2hw.tag_1734.re;
  assign rcache_line[6][198].status_reg.status = reg2hw.status_1734.q;//status_reg_t'(reg2hw.status_1734.q);
  assign rcache_line[6][198].status_reg.qe    = reg2hw.status_1734.qe;
  assign rcache_line[6][198].status_reg.re    = reg2hw.status_1734.re;


  assign rcache_line[6][199].tag_reg.tag      = reg2hw.tag_1735.q;
  assign rcache_line[6][199].tag_reg.qe       = reg2hw.tag_1735.qe;
  assign rcache_line[6][199].tag_reg.re       = reg2hw.tag_1735.re;
  assign rcache_line[6][199].status_reg.status = reg2hw.status_1735.q;//status_reg_t'(reg2hw.status_1735.q);
  assign rcache_line[6][199].status_reg.qe    = reg2hw.status_1735.qe;
  assign rcache_line[6][199].status_reg.re    = reg2hw.status_1735.re;


  assign rcache_line[6][200].tag_reg.tag      = reg2hw.tag_1736.q;
  assign rcache_line[6][200].tag_reg.qe       = reg2hw.tag_1736.qe;
  assign rcache_line[6][200].tag_reg.re       = reg2hw.tag_1736.re;
  assign rcache_line[6][200].status_reg.status = reg2hw.status_1736.q;//status_reg_t'(reg2hw.status_1736.q);
  assign rcache_line[6][200].status_reg.qe    = reg2hw.status_1736.qe;
  assign rcache_line[6][200].status_reg.re    = reg2hw.status_1736.re;


  assign rcache_line[6][201].tag_reg.tag      = reg2hw.tag_1737.q;
  assign rcache_line[6][201].tag_reg.qe       = reg2hw.tag_1737.qe;
  assign rcache_line[6][201].tag_reg.re       = reg2hw.tag_1737.re;
  assign rcache_line[6][201].status_reg.status = reg2hw.status_1737.q;//status_reg_t'(reg2hw.status_1737.q);
  assign rcache_line[6][201].status_reg.qe    = reg2hw.status_1737.qe;
  assign rcache_line[6][201].status_reg.re    = reg2hw.status_1737.re;


  assign rcache_line[6][202].tag_reg.tag      = reg2hw.tag_1738.q;
  assign rcache_line[6][202].tag_reg.qe       = reg2hw.tag_1738.qe;
  assign rcache_line[6][202].tag_reg.re       = reg2hw.tag_1738.re;
  assign rcache_line[6][202].status_reg.status = reg2hw.status_1738.q;//status_reg_t'(reg2hw.status_1738.q);
  assign rcache_line[6][202].status_reg.qe    = reg2hw.status_1738.qe;
  assign rcache_line[6][202].status_reg.re    = reg2hw.status_1738.re;


  assign rcache_line[6][203].tag_reg.tag      = reg2hw.tag_1739.q;
  assign rcache_line[6][203].tag_reg.qe       = reg2hw.tag_1739.qe;
  assign rcache_line[6][203].tag_reg.re       = reg2hw.tag_1739.re;
  assign rcache_line[6][203].status_reg.status = reg2hw.status_1739.q;//status_reg_t'(reg2hw.status_1739.q);
  assign rcache_line[6][203].status_reg.qe    = reg2hw.status_1739.qe;
  assign rcache_line[6][203].status_reg.re    = reg2hw.status_1739.re;


  assign rcache_line[6][204].tag_reg.tag      = reg2hw.tag_1740.q;
  assign rcache_line[6][204].tag_reg.qe       = reg2hw.tag_1740.qe;
  assign rcache_line[6][204].tag_reg.re       = reg2hw.tag_1740.re;
  assign rcache_line[6][204].status_reg.status = reg2hw.status_1740.q;//status_reg_t'(reg2hw.status_1740.q);
  assign rcache_line[6][204].status_reg.qe    = reg2hw.status_1740.qe;
  assign rcache_line[6][204].status_reg.re    = reg2hw.status_1740.re;


  assign rcache_line[6][205].tag_reg.tag      = reg2hw.tag_1741.q;
  assign rcache_line[6][205].tag_reg.qe       = reg2hw.tag_1741.qe;
  assign rcache_line[6][205].tag_reg.re       = reg2hw.tag_1741.re;
  assign rcache_line[6][205].status_reg.status = reg2hw.status_1741.q;//status_reg_t'(reg2hw.status_1741.q);
  assign rcache_line[6][205].status_reg.qe    = reg2hw.status_1741.qe;
  assign rcache_line[6][205].status_reg.re    = reg2hw.status_1741.re;


  assign rcache_line[6][206].tag_reg.tag      = reg2hw.tag_1742.q;
  assign rcache_line[6][206].tag_reg.qe       = reg2hw.tag_1742.qe;
  assign rcache_line[6][206].tag_reg.re       = reg2hw.tag_1742.re;
  assign rcache_line[6][206].status_reg.status = reg2hw.status_1742.q;//status_reg_t'(reg2hw.status_1742.q);
  assign rcache_line[6][206].status_reg.qe    = reg2hw.status_1742.qe;
  assign rcache_line[6][206].status_reg.re    = reg2hw.status_1742.re;


  assign rcache_line[6][207].tag_reg.tag      = reg2hw.tag_1743.q;
  assign rcache_line[6][207].tag_reg.qe       = reg2hw.tag_1743.qe;
  assign rcache_line[6][207].tag_reg.re       = reg2hw.tag_1743.re;
  assign rcache_line[6][207].status_reg.status = reg2hw.status_1743.q;//status_reg_t'(reg2hw.status_1743.q);
  assign rcache_line[6][207].status_reg.qe    = reg2hw.status_1743.qe;
  assign rcache_line[6][207].status_reg.re    = reg2hw.status_1743.re;


  assign rcache_line[6][208].tag_reg.tag      = reg2hw.tag_1744.q;
  assign rcache_line[6][208].tag_reg.qe       = reg2hw.tag_1744.qe;
  assign rcache_line[6][208].tag_reg.re       = reg2hw.tag_1744.re;
  assign rcache_line[6][208].status_reg.status = reg2hw.status_1744.q;//status_reg_t'(reg2hw.status_1744.q);
  assign rcache_line[6][208].status_reg.qe    = reg2hw.status_1744.qe;
  assign rcache_line[6][208].status_reg.re    = reg2hw.status_1744.re;


  assign rcache_line[6][209].tag_reg.tag      = reg2hw.tag_1745.q;
  assign rcache_line[6][209].tag_reg.qe       = reg2hw.tag_1745.qe;
  assign rcache_line[6][209].tag_reg.re       = reg2hw.tag_1745.re;
  assign rcache_line[6][209].status_reg.status = reg2hw.status_1745.q;//status_reg_t'(reg2hw.status_1745.q);
  assign rcache_line[6][209].status_reg.qe    = reg2hw.status_1745.qe;
  assign rcache_line[6][209].status_reg.re    = reg2hw.status_1745.re;


  assign rcache_line[6][210].tag_reg.tag      = reg2hw.tag_1746.q;
  assign rcache_line[6][210].tag_reg.qe       = reg2hw.tag_1746.qe;
  assign rcache_line[6][210].tag_reg.re       = reg2hw.tag_1746.re;
  assign rcache_line[6][210].status_reg.status = reg2hw.status_1746.q;//status_reg_t'(reg2hw.status_1746.q);
  assign rcache_line[6][210].status_reg.qe    = reg2hw.status_1746.qe;
  assign rcache_line[6][210].status_reg.re    = reg2hw.status_1746.re;


  assign rcache_line[6][211].tag_reg.tag      = reg2hw.tag_1747.q;
  assign rcache_line[6][211].tag_reg.qe       = reg2hw.tag_1747.qe;
  assign rcache_line[6][211].tag_reg.re       = reg2hw.tag_1747.re;
  assign rcache_line[6][211].status_reg.status = reg2hw.status_1747.q;//status_reg_t'(reg2hw.status_1747.q);
  assign rcache_line[6][211].status_reg.qe    = reg2hw.status_1747.qe;
  assign rcache_line[6][211].status_reg.re    = reg2hw.status_1747.re;


  assign rcache_line[6][212].tag_reg.tag      = reg2hw.tag_1748.q;
  assign rcache_line[6][212].tag_reg.qe       = reg2hw.tag_1748.qe;
  assign rcache_line[6][212].tag_reg.re       = reg2hw.tag_1748.re;
  assign rcache_line[6][212].status_reg.status = reg2hw.status_1748.q;//status_reg_t'(reg2hw.status_1748.q);
  assign rcache_line[6][212].status_reg.qe    = reg2hw.status_1748.qe;
  assign rcache_line[6][212].status_reg.re    = reg2hw.status_1748.re;


  assign rcache_line[6][213].tag_reg.tag      = reg2hw.tag_1749.q;
  assign rcache_line[6][213].tag_reg.qe       = reg2hw.tag_1749.qe;
  assign rcache_line[6][213].tag_reg.re       = reg2hw.tag_1749.re;
  assign rcache_line[6][213].status_reg.status = reg2hw.status_1749.q;//status_reg_t'(reg2hw.status_1749.q);
  assign rcache_line[6][213].status_reg.qe    = reg2hw.status_1749.qe;
  assign rcache_line[6][213].status_reg.re    = reg2hw.status_1749.re;


  assign rcache_line[6][214].tag_reg.tag      = reg2hw.tag_1750.q;
  assign rcache_line[6][214].tag_reg.qe       = reg2hw.tag_1750.qe;
  assign rcache_line[6][214].tag_reg.re       = reg2hw.tag_1750.re;
  assign rcache_line[6][214].status_reg.status = reg2hw.status_1750.q;//status_reg_t'(reg2hw.status_1750.q);
  assign rcache_line[6][214].status_reg.qe    = reg2hw.status_1750.qe;
  assign rcache_line[6][214].status_reg.re    = reg2hw.status_1750.re;


  assign rcache_line[6][215].tag_reg.tag      = reg2hw.tag_1751.q;
  assign rcache_line[6][215].tag_reg.qe       = reg2hw.tag_1751.qe;
  assign rcache_line[6][215].tag_reg.re       = reg2hw.tag_1751.re;
  assign rcache_line[6][215].status_reg.status = reg2hw.status_1751.q;//status_reg_t'(reg2hw.status_1751.q);
  assign rcache_line[6][215].status_reg.qe    = reg2hw.status_1751.qe;
  assign rcache_line[6][215].status_reg.re    = reg2hw.status_1751.re;


  assign rcache_line[6][216].tag_reg.tag      = reg2hw.tag_1752.q;
  assign rcache_line[6][216].tag_reg.qe       = reg2hw.tag_1752.qe;
  assign rcache_line[6][216].tag_reg.re       = reg2hw.tag_1752.re;
  assign rcache_line[6][216].status_reg.status = reg2hw.status_1752.q;//status_reg_t'(reg2hw.status_1752.q);
  assign rcache_line[6][216].status_reg.qe    = reg2hw.status_1752.qe;
  assign rcache_line[6][216].status_reg.re    = reg2hw.status_1752.re;


  assign rcache_line[6][217].tag_reg.tag      = reg2hw.tag_1753.q;
  assign rcache_line[6][217].tag_reg.qe       = reg2hw.tag_1753.qe;
  assign rcache_line[6][217].tag_reg.re       = reg2hw.tag_1753.re;
  assign rcache_line[6][217].status_reg.status = reg2hw.status_1753.q;//status_reg_t'(reg2hw.status_1753.q);
  assign rcache_line[6][217].status_reg.qe    = reg2hw.status_1753.qe;
  assign rcache_line[6][217].status_reg.re    = reg2hw.status_1753.re;


  assign rcache_line[6][218].tag_reg.tag      = reg2hw.tag_1754.q;
  assign rcache_line[6][218].tag_reg.qe       = reg2hw.tag_1754.qe;
  assign rcache_line[6][218].tag_reg.re       = reg2hw.tag_1754.re;
  assign rcache_line[6][218].status_reg.status = reg2hw.status_1754.q;//status_reg_t'(reg2hw.status_1754.q);
  assign rcache_line[6][218].status_reg.qe    = reg2hw.status_1754.qe;
  assign rcache_line[6][218].status_reg.re    = reg2hw.status_1754.re;


  assign rcache_line[6][219].tag_reg.tag      = reg2hw.tag_1755.q;
  assign rcache_line[6][219].tag_reg.qe       = reg2hw.tag_1755.qe;
  assign rcache_line[6][219].tag_reg.re       = reg2hw.tag_1755.re;
  assign rcache_line[6][219].status_reg.status = reg2hw.status_1755.q;//status_reg_t'(reg2hw.status_1755.q);
  assign rcache_line[6][219].status_reg.qe    = reg2hw.status_1755.qe;
  assign rcache_line[6][219].status_reg.re    = reg2hw.status_1755.re;


  assign rcache_line[6][220].tag_reg.tag      = reg2hw.tag_1756.q;
  assign rcache_line[6][220].tag_reg.qe       = reg2hw.tag_1756.qe;
  assign rcache_line[6][220].tag_reg.re       = reg2hw.tag_1756.re;
  assign rcache_line[6][220].status_reg.status = reg2hw.status_1756.q;//status_reg_t'(reg2hw.status_1756.q);
  assign rcache_line[6][220].status_reg.qe    = reg2hw.status_1756.qe;
  assign rcache_line[6][220].status_reg.re    = reg2hw.status_1756.re;


  assign rcache_line[6][221].tag_reg.tag      = reg2hw.tag_1757.q;
  assign rcache_line[6][221].tag_reg.qe       = reg2hw.tag_1757.qe;
  assign rcache_line[6][221].tag_reg.re       = reg2hw.tag_1757.re;
  assign rcache_line[6][221].status_reg.status = reg2hw.status_1757.q;//status_reg_t'(reg2hw.status_1757.q);
  assign rcache_line[6][221].status_reg.qe    = reg2hw.status_1757.qe;
  assign rcache_line[6][221].status_reg.re    = reg2hw.status_1757.re;


  assign rcache_line[6][222].tag_reg.tag      = reg2hw.tag_1758.q;
  assign rcache_line[6][222].tag_reg.qe       = reg2hw.tag_1758.qe;
  assign rcache_line[6][222].tag_reg.re       = reg2hw.tag_1758.re;
  assign rcache_line[6][222].status_reg.status = reg2hw.status_1758.q;//status_reg_t'(reg2hw.status_1758.q);
  assign rcache_line[6][222].status_reg.qe    = reg2hw.status_1758.qe;
  assign rcache_line[6][222].status_reg.re    = reg2hw.status_1758.re;


  assign rcache_line[6][223].tag_reg.tag      = reg2hw.tag_1759.q;
  assign rcache_line[6][223].tag_reg.qe       = reg2hw.tag_1759.qe;
  assign rcache_line[6][223].tag_reg.re       = reg2hw.tag_1759.re;
  assign rcache_line[6][223].status_reg.status = reg2hw.status_1759.q;//status_reg_t'(reg2hw.status_1759.q);
  assign rcache_line[6][223].status_reg.qe    = reg2hw.status_1759.qe;
  assign rcache_line[6][223].status_reg.re    = reg2hw.status_1759.re;


  assign rcache_line[6][224].tag_reg.tag      = reg2hw.tag_1760.q;
  assign rcache_line[6][224].tag_reg.qe       = reg2hw.tag_1760.qe;
  assign rcache_line[6][224].tag_reg.re       = reg2hw.tag_1760.re;
  assign rcache_line[6][224].status_reg.status = reg2hw.status_1760.q;//status_reg_t'(reg2hw.status_1760.q);
  assign rcache_line[6][224].status_reg.qe    = reg2hw.status_1760.qe;
  assign rcache_line[6][224].status_reg.re    = reg2hw.status_1760.re;


  assign rcache_line[6][225].tag_reg.tag      = reg2hw.tag_1761.q;
  assign rcache_line[6][225].tag_reg.qe       = reg2hw.tag_1761.qe;
  assign rcache_line[6][225].tag_reg.re       = reg2hw.tag_1761.re;
  assign rcache_line[6][225].status_reg.status = reg2hw.status_1761.q;//status_reg_t'(reg2hw.status_1761.q);
  assign rcache_line[6][225].status_reg.qe    = reg2hw.status_1761.qe;
  assign rcache_line[6][225].status_reg.re    = reg2hw.status_1761.re;


  assign rcache_line[6][226].tag_reg.tag      = reg2hw.tag_1762.q;
  assign rcache_line[6][226].tag_reg.qe       = reg2hw.tag_1762.qe;
  assign rcache_line[6][226].tag_reg.re       = reg2hw.tag_1762.re;
  assign rcache_line[6][226].status_reg.status = reg2hw.status_1762.q;//status_reg_t'(reg2hw.status_1762.q);
  assign rcache_line[6][226].status_reg.qe    = reg2hw.status_1762.qe;
  assign rcache_line[6][226].status_reg.re    = reg2hw.status_1762.re;


  assign rcache_line[6][227].tag_reg.tag      = reg2hw.tag_1763.q;
  assign rcache_line[6][227].tag_reg.qe       = reg2hw.tag_1763.qe;
  assign rcache_line[6][227].tag_reg.re       = reg2hw.tag_1763.re;
  assign rcache_line[6][227].status_reg.status = reg2hw.status_1763.q;//status_reg_t'(reg2hw.status_1763.q);
  assign rcache_line[6][227].status_reg.qe    = reg2hw.status_1763.qe;
  assign rcache_line[6][227].status_reg.re    = reg2hw.status_1763.re;


  assign rcache_line[6][228].tag_reg.tag      = reg2hw.tag_1764.q;
  assign rcache_line[6][228].tag_reg.qe       = reg2hw.tag_1764.qe;
  assign rcache_line[6][228].tag_reg.re       = reg2hw.tag_1764.re;
  assign rcache_line[6][228].status_reg.status = reg2hw.status_1764.q;//status_reg_t'(reg2hw.status_1764.q);
  assign rcache_line[6][228].status_reg.qe    = reg2hw.status_1764.qe;
  assign rcache_line[6][228].status_reg.re    = reg2hw.status_1764.re;


  assign rcache_line[6][229].tag_reg.tag      = reg2hw.tag_1765.q;
  assign rcache_line[6][229].tag_reg.qe       = reg2hw.tag_1765.qe;
  assign rcache_line[6][229].tag_reg.re       = reg2hw.tag_1765.re;
  assign rcache_line[6][229].status_reg.status = reg2hw.status_1765.q;//status_reg_t'(reg2hw.status_1765.q);
  assign rcache_line[6][229].status_reg.qe    = reg2hw.status_1765.qe;
  assign rcache_line[6][229].status_reg.re    = reg2hw.status_1765.re;


  assign rcache_line[6][230].tag_reg.tag      = reg2hw.tag_1766.q;
  assign rcache_line[6][230].tag_reg.qe       = reg2hw.tag_1766.qe;
  assign rcache_line[6][230].tag_reg.re       = reg2hw.tag_1766.re;
  assign rcache_line[6][230].status_reg.status = reg2hw.status_1766.q;//status_reg_t'(reg2hw.status_1766.q);
  assign rcache_line[6][230].status_reg.qe    = reg2hw.status_1766.qe;
  assign rcache_line[6][230].status_reg.re    = reg2hw.status_1766.re;


  assign rcache_line[6][231].tag_reg.tag      = reg2hw.tag_1767.q;
  assign rcache_line[6][231].tag_reg.qe       = reg2hw.tag_1767.qe;
  assign rcache_line[6][231].tag_reg.re       = reg2hw.tag_1767.re;
  assign rcache_line[6][231].status_reg.status = reg2hw.status_1767.q;//status_reg_t'(reg2hw.status_1767.q);
  assign rcache_line[6][231].status_reg.qe    = reg2hw.status_1767.qe;
  assign rcache_line[6][231].status_reg.re    = reg2hw.status_1767.re;


  assign rcache_line[6][232].tag_reg.tag      = reg2hw.tag_1768.q;
  assign rcache_line[6][232].tag_reg.qe       = reg2hw.tag_1768.qe;
  assign rcache_line[6][232].tag_reg.re       = reg2hw.tag_1768.re;
  assign rcache_line[6][232].status_reg.status = reg2hw.status_1768.q;//status_reg_t'(reg2hw.status_1768.q);
  assign rcache_line[6][232].status_reg.qe    = reg2hw.status_1768.qe;
  assign rcache_line[6][232].status_reg.re    = reg2hw.status_1768.re;


  assign rcache_line[6][233].tag_reg.tag      = reg2hw.tag_1769.q;
  assign rcache_line[6][233].tag_reg.qe       = reg2hw.tag_1769.qe;
  assign rcache_line[6][233].tag_reg.re       = reg2hw.tag_1769.re;
  assign rcache_line[6][233].status_reg.status = reg2hw.status_1769.q;//status_reg_t'(reg2hw.status_1769.q);
  assign rcache_line[6][233].status_reg.qe    = reg2hw.status_1769.qe;
  assign rcache_line[6][233].status_reg.re    = reg2hw.status_1769.re;


  assign rcache_line[6][234].tag_reg.tag      = reg2hw.tag_1770.q;
  assign rcache_line[6][234].tag_reg.qe       = reg2hw.tag_1770.qe;
  assign rcache_line[6][234].tag_reg.re       = reg2hw.tag_1770.re;
  assign rcache_line[6][234].status_reg.status = reg2hw.status_1770.q;//status_reg_t'(reg2hw.status_1770.q);
  assign rcache_line[6][234].status_reg.qe    = reg2hw.status_1770.qe;
  assign rcache_line[6][234].status_reg.re    = reg2hw.status_1770.re;


  assign rcache_line[6][235].tag_reg.tag      = reg2hw.tag_1771.q;
  assign rcache_line[6][235].tag_reg.qe       = reg2hw.tag_1771.qe;
  assign rcache_line[6][235].tag_reg.re       = reg2hw.tag_1771.re;
  assign rcache_line[6][235].status_reg.status = reg2hw.status_1771.q;//status_reg_t'(reg2hw.status_1771.q);
  assign rcache_line[6][235].status_reg.qe    = reg2hw.status_1771.qe;
  assign rcache_line[6][235].status_reg.re    = reg2hw.status_1771.re;


  assign rcache_line[6][236].tag_reg.tag      = reg2hw.tag_1772.q;
  assign rcache_line[6][236].tag_reg.qe       = reg2hw.tag_1772.qe;
  assign rcache_line[6][236].tag_reg.re       = reg2hw.tag_1772.re;
  assign rcache_line[6][236].status_reg.status = reg2hw.status_1772.q;//status_reg_t'(reg2hw.status_1772.q);
  assign rcache_line[6][236].status_reg.qe    = reg2hw.status_1772.qe;
  assign rcache_line[6][236].status_reg.re    = reg2hw.status_1772.re;


  assign rcache_line[6][237].tag_reg.tag      = reg2hw.tag_1773.q;
  assign rcache_line[6][237].tag_reg.qe       = reg2hw.tag_1773.qe;
  assign rcache_line[6][237].tag_reg.re       = reg2hw.tag_1773.re;
  assign rcache_line[6][237].status_reg.status = reg2hw.status_1773.q;//status_reg_t'(reg2hw.status_1773.q);
  assign rcache_line[6][237].status_reg.qe    = reg2hw.status_1773.qe;
  assign rcache_line[6][237].status_reg.re    = reg2hw.status_1773.re;


  assign rcache_line[6][238].tag_reg.tag      = reg2hw.tag_1774.q;
  assign rcache_line[6][238].tag_reg.qe       = reg2hw.tag_1774.qe;
  assign rcache_line[6][238].tag_reg.re       = reg2hw.tag_1774.re;
  assign rcache_line[6][238].status_reg.status = reg2hw.status_1774.q;//status_reg_t'(reg2hw.status_1774.q);
  assign rcache_line[6][238].status_reg.qe    = reg2hw.status_1774.qe;
  assign rcache_line[6][238].status_reg.re    = reg2hw.status_1774.re;


  assign rcache_line[6][239].tag_reg.tag      = reg2hw.tag_1775.q;
  assign rcache_line[6][239].tag_reg.qe       = reg2hw.tag_1775.qe;
  assign rcache_line[6][239].tag_reg.re       = reg2hw.tag_1775.re;
  assign rcache_line[6][239].status_reg.status = reg2hw.status_1775.q;//status_reg_t'(reg2hw.status_1775.q);
  assign rcache_line[6][239].status_reg.qe    = reg2hw.status_1775.qe;
  assign rcache_line[6][239].status_reg.re    = reg2hw.status_1775.re;


  assign rcache_line[6][240].tag_reg.tag      = reg2hw.tag_1776.q;
  assign rcache_line[6][240].tag_reg.qe       = reg2hw.tag_1776.qe;
  assign rcache_line[6][240].tag_reg.re       = reg2hw.tag_1776.re;
  assign rcache_line[6][240].status_reg.status = reg2hw.status_1776.q;//status_reg_t'(reg2hw.status_1776.q);
  assign rcache_line[6][240].status_reg.qe    = reg2hw.status_1776.qe;
  assign rcache_line[6][240].status_reg.re    = reg2hw.status_1776.re;


  assign rcache_line[6][241].tag_reg.tag      = reg2hw.tag_1777.q;
  assign rcache_line[6][241].tag_reg.qe       = reg2hw.tag_1777.qe;
  assign rcache_line[6][241].tag_reg.re       = reg2hw.tag_1777.re;
  assign rcache_line[6][241].status_reg.status = reg2hw.status_1777.q;//status_reg_t'(reg2hw.status_1777.q);
  assign rcache_line[6][241].status_reg.qe    = reg2hw.status_1777.qe;
  assign rcache_line[6][241].status_reg.re    = reg2hw.status_1777.re;


  assign rcache_line[6][242].tag_reg.tag      = reg2hw.tag_1778.q;
  assign rcache_line[6][242].tag_reg.qe       = reg2hw.tag_1778.qe;
  assign rcache_line[6][242].tag_reg.re       = reg2hw.tag_1778.re;
  assign rcache_line[6][242].status_reg.status = reg2hw.status_1778.q;//status_reg_t'(reg2hw.status_1778.q);
  assign rcache_line[6][242].status_reg.qe    = reg2hw.status_1778.qe;
  assign rcache_line[6][242].status_reg.re    = reg2hw.status_1778.re;


  assign rcache_line[6][243].tag_reg.tag      = reg2hw.tag_1779.q;
  assign rcache_line[6][243].tag_reg.qe       = reg2hw.tag_1779.qe;
  assign rcache_line[6][243].tag_reg.re       = reg2hw.tag_1779.re;
  assign rcache_line[6][243].status_reg.status = reg2hw.status_1779.q;//status_reg_t'(reg2hw.status_1779.q);
  assign rcache_line[6][243].status_reg.qe    = reg2hw.status_1779.qe;
  assign rcache_line[6][243].status_reg.re    = reg2hw.status_1779.re;


  assign rcache_line[6][244].tag_reg.tag      = reg2hw.tag_1780.q;
  assign rcache_line[6][244].tag_reg.qe       = reg2hw.tag_1780.qe;
  assign rcache_line[6][244].tag_reg.re       = reg2hw.tag_1780.re;
  assign rcache_line[6][244].status_reg.status = reg2hw.status_1780.q;//status_reg_t'(reg2hw.status_1780.q);
  assign rcache_line[6][244].status_reg.qe    = reg2hw.status_1780.qe;
  assign rcache_line[6][244].status_reg.re    = reg2hw.status_1780.re;


  assign rcache_line[6][245].tag_reg.tag      = reg2hw.tag_1781.q;
  assign rcache_line[6][245].tag_reg.qe       = reg2hw.tag_1781.qe;
  assign rcache_line[6][245].tag_reg.re       = reg2hw.tag_1781.re;
  assign rcache_line[6][245].status_reg.status = reg2hw.status_1781.q;//status_reg_t'(reg2hw.status_1781.q);
  assign rcache_line[6][245].status_reg.qe    = reg2hw.status_1781.qe;
  assign rcache_line[6][245].status_reg.re    = reg2hw.status_1781.re;


  assign rcache_line[6][246].tag_reg.tag      = reg2hw.tag_1782.q;
  assign rcache_line[6][246].tag_reg.qe       = reg2hw.tag_1782.qe;
  assign rcache_line[6][246].tag_reg.re       = reg2hw.tag_1782.re;
  assign rcache_line[6][246].status_reg.status = reg2hw.status_1782.q;//status_reg_t'(reg2hw.status_1782.q);
  assign rcache_line[6][246].status_reg.qe    = reg2hw.status_1782.qe;
  assign rcache_line[6][246].status_reg.re    = reg2hw.status_1782.re;


  assign rcache_line[6][247].tag_reg.tag      = reg2hw.tag_1783.q;
  assign rcache_line[6][247].tag_reg.qe       = reg2hw.tag_1783.qe;
  assign rcache_line[6][247].tag_reg.re       = reg2hw.tag_1783.re;
  assign rcache_line[6][247].status_reg.status = reg2hw.status_1783.q;//status_reg_t'(reg2hw.status_1783.q);
  assign rcache_line[6][247].status_reg.qe    = reg2hw.status_1783.qe;
  assign rcache_line[6][247].status_reg.re    = reg2hw.status_1783.re;


  assign rcache_line[6][248].tag_reg.tag      = reg2hw.tag_1784.q;
  assign rcache_line[6][248].tag_reg.qe       = reg2hw.tag_1784.qe;
  assign rcache_line[6][248].tag_reg.re       = reg2hw.tag_1784.re;
  assign rcache_line[6][248].status_reg.status = reg2hw.status_1784.q;//status_reg_t'(reg2hw.status_1784.q);
  assign rcache_line[6][248].status_reg.qe    = reg2hw.status_1784.qe;
  assign rcache_line[6][248].status_reg.re    = reg2hw.status_1784.re;


  assign rcache_line[6][249].tag_reg.tag      = reg2hw.tag_1785.q;
  assign rcache_line[6][249].tag_reg.qe       = reg2hw.tag_1785.qe;
  assign rcache_line[6][249].tag_reg.re       = reg2hw.tag_1785.re;
  assign rcache_line[6][249].status_reg.status = reg2hw.status_1785.q;//status_reg_t'(reg2hw.status_1785.q);
  assign rcache_line[6][249].status_reg.qe    = reg2hw.status_1785.qe;
  assign rcache_line[6][249].status_reg.re    = reg2hw.status_1785.re;


  assign rcache_line[6][250].tag_reg.tag      = reg2hw.tag_1786.q;
  assign rcache_line[6][250].tag_reg.qe       = reg2hw.tag_1786.qe;
  assign rcache_line[6][250].tag_reg.re       = reg2hw.tag_1786.re;
  assign rcache_line[6][250].status_reg.status = reg2hw.status_1786.q;//status_reg_t'(reg2hw.status_1786.q);
  assign rcache_line[6][250].status_reg.qe    = reg2hw.status_1786.qe;
  assign rcache_line[6][250].status_reg.re    = reg2hw.status_1786.re;


  assign rcache_line[6][251].tag_reg.tag      = reg2hw.tag_1787.q;
  assign rcache_line[6][251].tag_reg.qe       = reg2hw.tag_1787.qe;
  assign rcache_line[6][251].tag_reg.re       = reg2hw.tag_1787.re;
  assign rcache_line[6][251].status_reg.status = reg2hw.status_1787.q;//status_reg_t'(reg2hw.status_1787.q);
  assign rcache_line[6][251].status_reg.qe    = reg2hw.status_1787.qe;
  assign rcache_line[6][251].status_reg.re    = reg2hw.status_1787.re;


  assign rcache_line[6][252].tag_reg.tag      = reg2hw.tag_1788.q;
  assign rcache_line[6][252].tag_reg.qe       = reg2hw.tag_1788.qe;
  assign rcache_line[6][252].tag_reg.re       = reg2hw.tag_1788.re;
  assign rcache_line[6][252].status_reg.status = reg2hw.status_1788.q;//status_reg_t'(reg2hw.status_1788.q);
  assign rcache_line[6][252].status_reg.qe    = reg2hw.status_1788.qe;
  assign rcache_line[6][252].status_reg.re    = reg2hw.status_1788.re;


  assign rcache_line[6][253].tag_reg.tag      = reg2hw.tag_1789.q;
  assign rcache_line[6][253].tag_reg.qe       = reg2hw.tag_1789.qe;
  assign rcache_line[6][253].tag_reg.re       = reg2hw.tag_1789.re;
  assign rcache_line[6][253].status_reg.status = reg2hw.status_1789.q;//status_reg_t'(reg2hw.status_1789.q);
  assign rcache_line[6][253].status_reg.qe    = reg2hw.status_1789.qe;
  assign rcache_line[6][253].status_reg.re    = reg2hw.status_1789.re;


  assign rcache_line[6][254].tag_reg.tag      = reg2hw.tag_1790.q;
  assign rcache_line[6][254].tag_reg.qe       = reg2hw.tag_1790.qe;
  assign rcache_line[6][254].tag_reg.re       = reg2hw.tag_1790.re;
  assign rcache_line[6][254].status_reg.status = reg2hw.status_1790.q;//status_reg_t'(reg2hw.status_1790.q);
  assign rcache_line[6][254].status_reg.qe    = reg2hw.status_1790.qe;
  assign rcache_line[6][254].status_reg.re    = reg2hw.status_1790.re;


  assign rcache_line[6][255].tag_reg.tag      = reg2hw.tag_1791.q;
  assign rcache_line[6][255].tag_reg.qe       = reg2hw.tag_1791.qe;
  assign rcache_line[6][255].tag_reg.re       = reg2hw.tag_1791.re;
  assign rcache_line[6][255].status_reg.status = reg2hw.status_1791.q;//status_reg_t'(reg2hw.status_1791.q);
  assign rcache_line[6][255].status_reg.qe    = reg2hw.status_1791.qe;
  assign rcache_line[6][255].status_reg.re    = reg2hw.status_1791.re;


  assign rcache_line[7][0].tag_reg.tag      = reg2hw.tag_1792.q;
  assign rcache_line[7][0].tag_reg.qe       = reg2hw.tag_1792.qe;
  assign rcache_line[7][0].tag_reg.re       = reg2hw.tag_1792.re;
  assign rcache_line[7][0].status_reg.status = reg2hw.status_1792.q;//status_reg_t'(reg2hw.status_1792.q);
  assign rcache_line[7][0].status_reg.qe    = reg2hw.status_1792.qe;
  assign rcache_line[7][0].status_reg.re    = reg2hw.status_1792.re;


  assign rcache_line[7][1].tag_reg.tag      = reg2hw.tag_1793.q;
  assign rcache_line[7][1].tag_reg.qe       = reg2hw.tag_1793.qe;
  assign rcache_line[7][1].tag_reg.re       = reg2hw.tag_1793.re;
  assign rcache_line[7][1].status_reg.status = reg2hw.status_1793.q;//status_reg_t'(reg2hw.status_1793.q);
  assign rcache_line[7][1].status_reg.qe    = reg2hw.status_1793.qe;
  assign rcache_line[7][1].status_reg.re    = reg2hw.status_1793.re;


  assign rcache_line[7][2].tag_reg.tag      = reg2hw.tag_1794.q;
  assign rcache_line[7][2].tag_reg.qe       = reg2hw.tag_1794.qe;
  assign rcache_line[7][2].tag_reg.re       = reg2hw.tag_1794.re;
  assign rcache_line[7][2].status_reg.status = reg2hw.status_1794.q;//status_reg_t'(reg2hw.status_1794.q);
  assign rcache_line[7][2].status_reg.qe    = reg2hw.status_1794.qe;
  assign rcache_line[7][2].status_reg.re    = reg2hw.status_1794.re;


  assign rcache_line[7][3].tag_reg.tag      = reg2hw.tag_1795.q;
  assign rcache_line[7][3].tag_reg.qe       = reg2hw.tag_1795.qe;
  assign rcache_line[7][3].tag_reg.re       = reg2hw.tag_1795.re;
  assign rcache_line[7][3].status_reg.status = reg2hw.status_1795.q;//status_reg_t'(reg2hw.status_1795.q);
  assign rcache_line[7][3].status_reg.qe    = reg2hw.status_1795.qe;
  assign rcache_line[7][3].status_reg.re    = reg2hw.status_1795.re;


  assign rcache_line[7][4].tag_reg.tag      = reg2hw.tag_1796.q;
  assign rcache_line[7][4].tag_reg.qe       = reg2hw.tag_1796.qe;
  assign rcache_line[7][4].tag_reg.re       = reg2hw.tag_1796.re;
  assign rcache_line[7][4].status_reg.status = reg2hw.status_1796.q;//status_reg_t'(reg2hw.status_1796.q);
  assign rcache_line[7][4].status_reg.qe    = reg2hw.status_1796.qe;
  assign rcache_line[7][4].status_reg.re    = reg2hw.status_1796.re;


  assign rcache_line[7][5].tag_reg.tag      = reg2hw.tag_1797.q;
  assign rcache_line[7][5].tag_reg.qe       = reg2hw.tag_1797.qe;
  assign rcache_line[7][5].tag_reg.re       = reg2hw.tag_1797.re;
  assign rcache_line[7][5].status_reg.status = reg2hw.status_1797.q;//status_reg_t'(reg2hw.status_1797.q);
  assign rcache_line[7][5].status_reg.qe    = reg2hw.status_1797.qe;
  assign rcache_line[7][5].status_reg.re    = reg2hw.status_1797.re;


  assign rcache_line[7][6].tag_reg.tag      = reg2hw.tag_1798.q;
  assign rcache_line[7][6].tag_reg.qe       = reg2hw.tag_1798.qe;
  assign rcache_line[7][6].tag_reg.re       = reg2hw.tag_1798.re;
  assign rcache_line[7][6].status_reg.status = reg2hw.status_1798.q;//status_reg_t'(reg2hw.status_1798.q);
  assign rcache_line[7][6].status_reg.qe    = reg2hw.status_1798.qe;
  assign rcache_line[7][6].status_reg.re    = reg2hw.status_1798.re;


  assign rcache_line[7][7].tag_reg.tag      = reg2hw.tag_1799.q;
  assign rcache_line[7][7].tag_reg.qe       = reg2hw.tag_1799.qe;
  assign rcache_line[7][7].tag_reg.re       = reg2hw.tag_1799.re;
  assign rcache_line[7][7].status_reg.status = reg2hw.status_1799.q;//status_reg_t'(reg2hw.status_1799.q);
  assign rcache_line[7][7].status_reg.qe    = reg2hw.status_1799.qe;
  assign rcache_line[7][7].status_reg.re    = reg2hw.status_1799.re;


  assign rcache_line[7][8].tag_reg.tag      = reg2hw.tag_1800.q;
  assign rcache_line[7][8].tag_reg.qe       = reg2hw.tag_1800.qe;
  assign rcache_line[7][8].tag_reg.re       = reg2hw.tag_1800.re;
  assign rcache_line[7][8].status_reg.status = reg2hw.status_1800.q;//status_reg_t'(reg2hw.status_1800.q);
  assign rcache_line[7][8].status_reg.qe    = reg2hw.status_1800.qe;
  assign rcache_line[7][8].status_reg.re    = reg2hw.status_1800.re;


  assign rcache_line[7][9].tag_reg.tag      = reg2hw.tag_1801.q;
  assign rcache_line[7][9].tag_reg.qe       = reg2hw.tag_1801.qe;
  assign rcache_line[7][9].tag_reg.re       = reg2hw.tag_1801.re;
  assign rcache_line[7][9].status_reg.status = reg2hw.status_1801.q;//status_reg_t'(reg2hw.status_1801.q);
  assign rcache_line[7][9].status_reg.qe    = reg2hw.status_1801.qe;
  assign rcache_line[7][9].status_reg.re    = reg2hw.status_1801.re;


  assign rcache_line[7][10].tag_reg.tag      = reg2hw.tag_1802.q;
  assign rcache_line[7][10].tag_reg.qe       = reg2hw.tag_1802.qe;
  assign rcache_line[7][10].tag_reg.re       = reg2hw.tag_1802.re;
  assign rcache_line[7][10].status_reg.status = reg2hw.status_1802.q;//status_reg_t'(reg2hw.status_1802.q);
  assign rcache_line[7][10].status_reg.qe    = reg2hw.status_1802.qe;
  assign rcache_line[7][10].status_reg.re    = reg2hw.status_1802.re;


  assign rcache_line[7][11].tag_reg.tag      = reg2hw.tag_1803.q;
  assign rcache_line[7][11].tag_reg.qe       = reg2hw.tag_1803.qe;
  assign rcache_line[7][11].tag_reg.re       = reg2hw.tag_1803.re;
  assign rcache_line[7][11].status_reg.status = reg2hw.status_1803.q;//status_reg_t'(reg2hw.status_1803.q);
  assign rcache_line[7][11].status_reg.qe    = reg2hw.status_1803.qe;
  assign rcache_line[7][11].status_reg.re    = reg2hw.status_1803.re;


  assign rcache_line[7][12].tag_reg.tag      = reg2hw.tag_1804.q;
  assign rcache_line[7][12].tag_reg.qe       = reg2hw.tag_1804.qe;
  assign rcache_line[7][12].tag_reg.re       = reg2hw.tag_1804.re;
  assign rcache_line[7][12].status_reg.status = reg2hw.status_1804.q;//status_reg_t'(reg2hw.status_1804.q);
  assign rcache_line[7][12].status_reg.qe    = reg2hw.status_1804.qe;
  assign rcache_line[7][12].status_reg.re    = reg2hw.status_1804.re;


  assign rcache_line[7][13].tag_reg.tag      = reg2hw.tag_1805.q;
  assign rcache_line[7][13].tag_reg.qe       = reg2hw.tag_1805.qe;
  assign rcache_line[7][13].tag_reg.re       = reg2hw.tag_1805.re;
  assign rcache_line[7][13].status_reg.status = reg2hw.status_1805.q;//status_reg_t'(reg2hw.status_1805.q);
  assign rcache_line[7][13].status_reg.qe    = reg2hw.status_1805.qe;
  assign rcache_line[7][13].status_reg.re    = reg2hw.status_1805.re;


  assign rcache_line[7][14].tag_reg.tag      = reg2hw.tag_1806.q;
  assign rcache_line[7][14].tag_reg.qe       = reg2hw.tag_1806.qe;
  assign rcache_line[7][14].tag_reg.re       = reg2hw.tag_1806.re;
  assign rcache_line[7][14].status_reg.status = reg2hw.status_1806.q;//status_reg_t'(reg2hw.status_1806.q);
  assign rcache_line[7][14].status_reg.qe    = reg2hw.status_1806.qe;
  assign rcache_line[7][14].status_reg.re    = reg2hw.status_1806.re;


  assign rcache_line[7][15].tag_reg.tag      = reg2hw.tag_1807.q;
  assign rcache_line[7][15].tag_reg.qe       = reg2hw.tag_1807.qe;
  assign rcache_line[7][15].tag_reg.re       = reg2hw.tag_1807.re;
  assign rcache_line[7][15].status_reg.status = reg2hw.status_1807.q;//status_reg_t'(reg2hw.status_1807.q);
  assign rcache_line[7][15].status_reg.qe    = reg2hw.status_1807.qe;
  assign rcache_line[7][15].status_reg.re    = reg2hw.status_1807.re;


  assign rcache_line[7][16].tag_reg.tag      = reg2hw.tag_1808.q;
  assign rcache_line[7][16].tag_reg.qe       = reg2hw.tag_1808.qe;
  assign rcache_line[7][16].tag_reg.re       = reg2hw.tag_1808.re;
  assign rcache_line[7][16].status_reg.status = reg2hw.status_1808.q;//status_reg_t'(reg2hw.status_1808.q);
  assign rcache_line[7][16].status_reg.qe    = reg2hw.status_1808.qe;
  assign rcache_line[7][16].status_reg.re    = reg2hw.status_1808.re;


  assign rcache_line[7][17].tag_reg.tag      = reg2hw.tag_1809.q;
  assign rcache_line[7][17].tag_reg.qe       = reg2hw.tag_1809.qe;
  assign rcache_line[7][17].tag_reg.re       = reg2hw.tag_1809.re;
  assign rcache_line[7][17].status_reg.status = reg2hw.status_1809.q;//status_reg_t'(reg2hw.status_1809.q);
  assign rcache_line[7][17].status_reg.qe    = reg2hw.status_1809.qe;
  assign rcache_line[7][17].status_reg.re    = reg2hw.status_1809.re;


  assign rcache_line[7][18].tag_reg.tag      = reg2hw.tag_1810.q;
  assign rcache_line[7][18].tag_reg.qe       = reg2hw.tag_1810.qe;
  assign rcache_line[7][18].tag_reg.re       = reg2hw.tag_1810.re;
  assign rcache_line[7][18].status_reg.status = reg2hw.status_1810.q;//status_reg_t'(reg2hw.status_1810.q);
  assign rcache_line[7][18].status_reg.qe    = reg2hw.status_1810.qe;
  assign rcache_line[7][18].status_reg.re    = reg2hw.status_1810.re;


  assign rcache_line[7][19].tag_reg.tag      = reg2hw.tag_1811.q;
  assign rcache_line[7][19].tag_reg.qe       = reg2hw.tag_1811.qe;
  assign rcache_line[7][19].tag_reg.re       = reg2hw.tag_1811.re;
  assign rcache_line[7][19].status_reg.status = reg2hw.status_1811.q;//status_reg_t'(reg2hw.status_1811.q);
  assign rcache_line[7][19].status_reg.qe    = reg2hw.status_1811.qe;
  assign rcache_line[7][19].status_reg.re    = reg2hw.status_1811.re;


  assign rcache_line[7][20].tag_reg.tag      = reg2hw.tag_1812.q;
  assign rcache_line[7][20].tag_reg.qe       = reg2hw.tag_1812.qe;
  assign rcache_line[7][20].tag_reg.re       = reg2hw.tag_1812.re;
  assign rcache_line[7][20].status_reg.status = reg2hw.status_1812.q;//status_reg_t'(reg2hw.status_1812.q);
  assign rcache_line[7][20].status_reg.qe    = reg2hw.status_1812.qe;
  assign rcache_line[7][20].status_reg.re    = reg2hw.status_1812.re;


  assign rcache_line[7][21].tag_reg.tag      = reg2hw.tag_1813.q;
  assign rcache_line[7][21].tag_reg.qe       = reg2hw.tag_1813.qe;
  assign rcache_line[7][21].tag_reg.re       = reg2hw.tag_1813.re;
  assign rcache_line[7][21].status_reg.status = reg2hw.status_1813.q;//status_reg_t'(reg2hw.status_1813.q);
  assign rcache_line[7][21].status_reg.qe    = reg2hw.status_1813.qe;
  assign rcache_line[7][21].status_reg.re    = reg2hw.status_1813.re;


  assign rcache_line[7][22].tag_reg.tag      = reg2hw.tag_1814.q;
  assign rcache_line[7][22].tag_reg.qe       = reg2hw.tag_1814.qe;
  assign rcache_line[7][22].tag_reg.re       = reg2hw.tag_1814.re;
  assign rcache_line[7][22].status_reg.status = reg2hw.status_1814.q;//status_reg_t'(reg2hw.status_1814.q);
  assign rcache_line[7][22].status_reg.qe    = reg2hw.status_1814.qe;
  assign rcache_line[7][22].status_reg.re    = reg2hw.status_1814.re;


  assign rcache_line[7][23].tag_reg.tag      = reg2hw.tag_1815.q;
  assign rcache_line[7][23].tag_reg.qe       = reg2hw.tag_1815.qe;
  assign rcache_line[7][23].tag_reg.re       = reg2hw.tag_1815.re;
  assign rcache_line[7][23].status_reg.status = reg2hw.status_1815.q;//status_reg_t'(reg2hw.status_1815.q);
  assign rcache_line[7][23].status_reg.qe    = reg2hw.status_1815.qe;
  assign rcache_line[7][23].status_reg.re    = reg2hw.status_1815.re;


  assign rcache_line[7][24].tag_reg.tag      = reg2hw.tag_1816.q;
  assign rcache_line[7][24].tag_reg.qe       = reg2hw.tag_1816.qe;
  assign rcache_line[7][24].tag_reg.re       = reg2hw.tag_1816.re;
  assign rcache_line[7][24].status_reg.status = reg2hw.status_1816.q;//status_reg_t'(reg2hw.status_1816.q);
  assign rcache_line[7][24].status_reg.qe    = reg2hw.status_1816.qe;
  assign rcache_line[7][24].status_reg.re    = reg2hw.status_1816.re;


  assign rcache_line[7][25].tag_reg.tag      = reg2hw.tag_1817.q;
  assign rcache_line[7][25].tag_reg.qe       = reg2hw.tag_1817.qe;
  assign rcache_line[7][25].tag_reg.re       = reg2hw.tag_1817.re;
  assign rcache_line[7][25].status_reg.status = reg2hw.status_1817.q;//status_reg_t'(reg2hw.status_1817.q);
  assign rcache_line[7][25].status_reg.qe    = reg2hw.status_1817.qe;
  assign rcache_line[7][25].status_reg.re    = reg2hw.status_1817.re;


  assign rcache_line[7][26].tag_reg.tag      = reg2hw.tag_1818.q;
  assign rcache_line[7][26].tag_reg.qe       = reg2hw.tag_1818.qe;
  assign rcache_line[7][26].tag_reg.re       = reg2hw.tag_1818.re;
  assign rcache_line[7][26].status_reg.status = reg2hw.status_1818.q;//status_reg_t'(reg2hw.status_1818.q);
  assign rcache_line[7][26].status_reg.qe    = reg2hw.status_1818.qe;
  assign rcache_line[7][26].status_reg.re    = reg2hw.status_1818.re;


  assign rcache_line[7][27].tag_reg.tag      = reg2hw.tag_1819.q;
  assign rcache_line[7][27].tag_reg.qe       = reg2hw.tag_1819.qe;
  assign rcache_line[7][27].tag_reg.re       = reg2hw.tag_1819.re;
  assign rcache_line[7][27].status_reg.status = reg2hw.status_1819.q;//status_reg_t'(reg2hw.status_1819.q);
  assign rcache_line[7][27].status_reg.qe    = reg2hw.status_1819.qe;
  assign rcache_line[7][27].status_reg.re    = reg2hw.status_1819.re;


  assign rcache_line[7][28].tag_reg.tag      = reg2hw.tag_1820.q;
  assign rcache_line[7][28].tag_reg.qe       = reg2hw.tag_1820.qe;
  assign rcache_line[7][28].tag_reg.re       = reg2hw.tag_1820.re;
  assign rcache_line[7][28].status_reg.status = reg2hw.status_1820.q;//status_reg_t'(reg2hw.status_1820.q);
  assign rcache_line[7][28].status_reg.qe    = reg2hw.status_1820.qe;
  assign rcache_line[7][28].status_reg.re    = reg2hw.status_1820.re;


  assign rcache_line[7][29].tag_reg.tag      = reg2hw.tag_1821.q;
  assign rcache_line[7][29].tag_reg.qe       = reg2hw.tag_1821.qe;
  assign rcache_line[7][29].tag_reg.re       = reg2hw.tag_1821.re;
  assign rcache_line[7][29].status_reg.status = reg2hw.status_1821.q;//status_reg_t'(reg2hw.status_1821.q);
  assign rcache_line[7][29].status_reg.qe    = reg2hw.status_1821.qe;
  assign rcache_line[7][29].status_reg.re    = reg2hw.status_1821.re;


  assign rcache_line[7][30].tag_reg.tag      = reg2hw.tag_1822.q;
  assign rcache_line[7][30].tag_reg.qe       = reg2hw.tag_1822.qe;
  assign rcache_line[7][30].tag_reg.re       = reg2hw.tag_1822.re;
  assign rcache_line[7][30].status_reg.status = reg2hw.status_1822.q;//status_reg_t'(reg2hw.status_1822.q);
  assign rcache_line[7][30].status_reg.qe    = reg2hw.status_1822.qe;
  assign rcache_line[7][30].status_reg.re    = reg2hw.status_1822.re;


  assign rcache_line[7][31].tag_reg.tag      = reg2hw.tag_1823.q;
  assign rcache_line[7][31].tag_reg.qe       = reg2hw.tag_1823.qe;
  assign rcache_line[7][31].tag_reg.re       = reg2hw.tag_1823.re;
  assign rcache_line[7][31].status_reg.status = reg2hw.status_1823.q;//status_reg_t'(reg2hw.status_1823.q);
  assign rcache_line[7][31].status_reg.qe    = reg2hw.status_1823.qe;
  assign rcache_line[7][31].status_reg.re    = reg2hw.status_1823.re;


  assign rcache_line[7][32].tag_reg.tag      = reg2hw.tag_1824.q;
  assign rcache_line[7][32].tag_reg.qe       = reg2hw.tag_1824.qe;
  assign rcache_line[7][32].tag_reg.re       = reg2hw.tag_1824.re;
  assign rcache_line[7][32].status_reg.status = reg2hw.status_1824.q;//status_reg_t'(reg2hw.status_1824.q);
  assign rcache_line[7][32].status_reg.qe    = reg2hw.status_1824.qe;
  assign rcache_line[7][32].status_reg.re    = reg2hw.status_1824.re;


  assign rcache_line[7][33].tag_reg.tag      = reg2hw.tag_1825.q;
  assign rcache_line[7][33].tag_reg.qe       = reg2hw.tag_1825.qe;
  assign rcache_line[7][33].tag_reg.re       = reg2hw.tag_1825.re;
  assign rcache_line[7][33].status_reg.status = reg2hw.status_1825.q;//status_reg_t'(reg2hw.status_1825.q);
  assign rcache_line[7][33].status_reg.qe    = reg2hw.status_1825.qe;
  assign rcache_line[7][33].status_reg.re    = reg2hw.status_1825.re;


  assign rcache_line[7][34].tag_reg.tag      = reg2hw.tag_1826.q;
  assign rcache_line[7][34].tag_reg.qe       = reg2hw.tag_1826.qe;
  assign rcache_line[7][34].tag_reg.re       = reg2hw.tag_1826.re;
  assign rcache_line[7][34].status_reg.status = reg2hw.status_1826.q;//status_reg_t'(reg2hw.status_1826.q);
  assign rcache_line[7][34].status_reg.qe    = reg2hw.status_1826.qe;
  assign rcache_line[7][34].status_reg.re    = reg2hw.status_1826.re;


  assign rcache_line[7][35].tag_reg.tag      = reg2hw.tag_1827.q;
  assign rcache_line[7][35].tag_reg.qe       = reg2hw.tag_1827.qe;
  assign rcache_line[7][35].tag_reg.re       = reg2hw.tag_1827.re;
  assign rcache_line[7][35].status_reg.status = reg2hw.status_1827.q;//status_reg_t'(reg2hw.status_1827.q);
  assign rcache_line[7][35].status_reg.qe    = reg2hw.status_1827.qe;
  assign rcache_line[7][35].status_reg.re    = reg2hw.status_1827.re;


  assign rcache_line[7][36].tag_reg.tag      = reg2hw.tag_1828.q;
  assign rcache_line[7][36].tag_reg.qe       = reg2hw.tag_1828.qe;
  assign rcache_line[7][36].tag_reg.re       = reg2hw.tag_1828.re;
  assign rcache_line[7][36].status_reg.status = reg2hw.status_1828.q;//status_reg_t'(reg2hw.status_1828.q);
  assign rcache_line[7][36].status_reg.qe    = reg2hw.status_1828.qe;
  assign rcache_line[7][36].status_reg.re    = reg2hw.status_1828.re;


  assign rcache_line[7][37].tag_reg.tag      = reg2hw.tag_1829.q;
  assign rcache_line[7][37].tag_reg.qe       = reg2hw.tag_1829.qe;
  assign rcache_line[7][37].tag_reg.re       = reg2hw.tag_1829.re;
  assign rcache_line[7][37].status_reg.status = reg2hw.status_1829.q;//status_reg_t'(reg2hw.status_1829.q);
  assign rcache_line[7][37].status_reg.qe    = reg2hw.status_1829.qe;
  assign rcache_line[7][37].status_reg.re    = reg2hw.status_1829.re;


  assign rcache_line[7][38].tag_reg.tag      = reg2hw.tag_1830.q;
  assign rcache_line[7][38].tag_reg.qe       = reg2hw.tag_1830.qe;
  assign rcache_line[7][38].tag_reg.re       = reg2hw.tag_1830.re;
  assign rcache_line[7][38].status_reg.status = reg2hw.status_1830.q;//status_reg_t'(reg2hw.status_1830.q);
  assign rcache_line[7][38].status_reg.qe    = reg2hw.status_1830.qe;
  assign rcache_line[7][38].status_reg.re    = reg2hw.status_1830.re;


  assign rcache_line[7][39].tag_reg.tag      = reg2hw.tag_1831.q;
  assign rcache_line[7][39].tag_reg.qe       = reg2hw.tag_1831.qe;
  assign rcache_line[7][39].tag_reg.re       = reg2hw.tag_1831.re;
  assign rcache_line[7][39].status_reg.status = reg2hw.status_1831.q;//status_reg_t'(reg2hw.status_1831.q);
  assign rcache_line[7][39].status_reg.qe    = reg2hw.status_1831.qe;
  assign rcache_line[7][39].status_reg.re    = reg2hw.status_1831.re;


  assign rcache_line[7][40].tag_reg.tag      = reg2hw.tag_1832.q;
  assign rcache_line[7][40].tag_reg.qe       = reg2hw.tag_1832.qe;
  assign rcache_line[7][40].tag_reg.re       = reg2hw.tag_1832.re;
  assign rcache_line[7][40].status_reg.status = reg2hw.status_1832.q;//status_reg_t'(reg2hw.status_1832.q);
  assign rcache_line[7][40].status_reg.qe    = reg2hw.status_1832.qe;
  assign rcache_line[7][40].status_reg.re    = reg2hw.status_1832.re;


  assign rcache_line[7][41].tag_reg.tag      = reg2hw.tag_1833.q;
  assign rcache_line[7][41].tag_reg.qe       = reg2hw.tag_1833.qe;
  assign rcache_line[7][41].tag_reg.re       = reg2hw.tag_1833.re;
  assign rcache_line[7][41].status_reg.status = reg2hw.status_1833.q;//status_reg_t'(reg2hw.status_1833.q);
  assign rcache_line[7][41].status_reg.qe    = reg2hw.status_1833.qe;
  assign rcache_line[7][41].status_reg.re    = reg2hw.status_1833.re;


  assign rcache_line[7][42].tag_reg.tag      = reg2hw.tag_1834.q;
  assign rcache_line[7][42].tag_reg.qe       = reg2hw.tag_1834.qe;
  assign rcache_line[7][42].tag_reg.re       = reg2hw.tag_1834.re;
  assign rcache_line[7][42].status_reg.status = reg2hw.status_1834.q;//status_reg_t'(reg2hw.status_1834.q);
  assign rcache_line[7][42].status_reg.qe    = reg2hw.status_1834.qe;
  assign rcache_line[7][42].status_reg.re    = reg2hw.status_1834.re;


  assign rcache_line[7][43].tag_reg.tag      = reg2hw.tag_1835.q;
  assign rcache_line[7][43].tag_reg.qe       = reg2hw.tag_1835.qe;
  assign rcache_line[7][43].tag_reg.re       = reg2hw.tag_1835.re;
  assign rcache_line[7][43].status_reg.status = reg2hw.status_1835.q;//status_reg_t'(reg2hw.status_1835.q);
  assign rcache_line[7][43].status_reg.qe    = reg2hw.status_1835.qe;
  assign rcache_line[7][43].status_reg.re    = reg2hw.status_1835.re;


  assign rcache_line[7][44].tag_reg.tag      = reg2hw.tag_1836.q;
  assign rcache_line[7][44].tag_reg.qe       = reg2hw.tag_1836.qe;
  assign rcache_line[7][44].tag_reg.re       = reg2hw.tag_1836.re;
  assign rcache_line[7][44].status_reg.status = reg2hw.status_1836.q;//status_reg_t'(reg2hw.status_1836.q);
  assign rcache_line[7][44].status_reg.qe    = reg2hw.status_1836.qe;
  assign rcache_line[7][44].status_reg.re    = reg2hw.status_1836.re;


  assign rcache_line[7][45].tag_reg.tag      = reg2hw.tag_1837.q;
  assign rcache_line[7][45].tag_reg.qe       = reg2hw.tag_1837.qe;
  assign rcache_line[7][45].tag_reg.re       = reg2hw.tag_1837.re;
  assign rcache_line[7][45].status_reg.status = reg2hw.status_1837.q;//status_reg_t'(reg2hw.status_1837.q);
  assign rcache_line[7][45].status_reg.qe    = reg2hw.status_1837.qe;
  assign rcache_line[7][45].status_reg.re    = reg2hw.status_1837.re;


  assign rcache_line[7][46].tag_reg.tag      = reg2hw.tag_1838.q;
  assign rcache_line[7][46].tag_reg.qe       = reg2hw.tag_1838.qe;
  assign rcache_line[7][46].tag_reg.re       = reg2hw.tag_1838.re;
  assign rcache_line[7][46].status_reg.status = reg2hw.status_1838.q;//status_reg_t'(reg2hw.status_1838.q);
  assign rcache_line[7][46].status_reg.qe    = reg2hw.status_1838.qe;
  assign rcache_line[7][46].status_reg.re    = reg2hw.status_1838.re;


  assign rcache_line[7][47].tag_reg.tag      = reg2hw.tag_1839.q;
  assign rcache_line[7][47].tag_reg.qe       = reg2hw.tag_1839.qe;
  assign rcache_line[7][47].tag_reg.re       = reg2hw.tag_1839.re;
  assign rcache_line[7][47].status_reg.status = reg2hw.status_1839.q;//status_reg_t'(reg2hw.status_1839.q);
  assign rcache_line[7][47].status_reg.qe    = reg2hw.status_1839.qe;
  assign rcache_line[7][47].status_reg.re    = reg2hw.status_1839.re;


  assign rcache_line[7][48].tag_reg.tag      = reg2hw.tag_1840.q;
  assign rcache_line[7][48].tag_reg.qe       = reg2hw.tag_1840.qe;
  assign rcache_line[7][48].tag_reg.re       = reg2hw.tag_1840.re;
  assign rcache_line[7][48].status_reg.status = reg2hw.status_1840.q;//status_reg_t'(reg2hw.status_1840.q);
  assign rcache_line[7][48].status_reg.qe    = reg2hw.status_1840.qe;
  assign rcache_line[7][48].status_reg.re    = reg2hw.status_1840.re;


  assign rcache_line[7][49].tag_reg.tag      = reg2hw.tag_1841.q;
  assign rcache_line[7][49].tag_reg.qe       = reg2hw.tag_1841.qe;
  assign rcache_line[7][49].tag_reg.re       = reg2hw.tag_1841.re;
  assign rcache_line[7][49].status_reg.status = reg2hw.status_1841.q;//status_reg_t'(reg2hw.status_1841.q);
  assign rcache_line[7][49].status_reg.qe    = reg2hw.status_1841.qe;
  assign rcache_line[7][49].status_reg.re    = reg2hw.status_1841.re;


  assign rcache_line[7][50].tag_reg.tag      = reg2hw.tag_1842.q;
  assign rcache_line[7][50].tag_reg.qe       = reg2hw.tag_1842.qe;
  assign rcache_line[7][50].tag_reg.re       = reg2hw.tag_1842.re;
  assign rcache_line[7][50].status_reg.status = reg2hw.status_1842.q;//status_reg_t'(reg2hw.status_1842.q);
  assign rcache_line[7][50].status_reg.qe    = reg2hw.status_1842.qe;
  assign rcache_line[7][50].status_reg.re    = reg2hw.status_1842.re;


  assign rcache_line[7][51].tag_reg.tag      = reg2hw.tag_1843.q;
  assign rcache_line[7][51].tag_reg.qe       = reg2hw.tag_1843.qe;
  assign rcache_line[7][51].tag_reg.re       = reg2hw.tag_1843.re;
  assign rcache_line[7][51].status_reg.status = reg2hw.status_1843.q;//status_reg_t'(reg2hw.status_1843.q);
  assign rcache_line[7][51].status_reg.qe    = reg2hw.status_1843.qe;
  assign rcache_line[7][51].status_reg.re    = reg2hw.status_1843.re;


  assign rcache_line[7][52].tag_reg.tag      = reg2hw.tag_1844.q;
  assign rcache_line[7][52].tag_reg.qe       = reg2hw.tag_1844.qe;
  assign rcache_line[7][52].tag_reg.re       = reg2hw.tag_1844.re;
  assign rcache_line[7][52].status_reg.status = reg2hw.status_1844.q;//status_reg_t'(reg2hw.status_1844.q);
  assign rcache_line[7][52].status_reg.qe    = reg2hw.status_1844.qe;
  assign rcache_line[7][52].status_reg.re    = reg2hw.status_1844.re;


  assign rcache_line[7][53].tag_reg.tag      = reg2hw.tag_1845.q;
  assign rcache_line[7][53].tag_reg.qe       = reg2hw.tag_1845.qe;
  assign rcache_line[7][53].tag_reg.re       = reg2hw.tag_1845.re;
  assign rcache_line[7][53].status_reg.status = reg2hw.status_1845.q;//status_reg_t'(reg2hw.status_1845.q);
  assign rcache_line[7][53].status_reg.qe    = reg2hw.status_1845.qe;
  assign rcache_line[7][53].status_reg.re    = reg2hw.status_1845.re;


  assign rcache_line[7][54].tag_reg.tag      = reg2hw.tag_1846.q;
  assign rcache_line[7][54].tag_reg.qe       = reg2hw.tag_1846.qe;
  assign rcache_line[7][54].tag_reg.re       = reg2hw.tag_1846.re;
  assign rcache_line[7][54].status_reg.status = reg2hw.status_1846.q;//status_reg_t'(reg2hw.status_1846.q);
  assign rcache_line[7][54].status_reg.qe    = reg2hw.status_1846.qe;
  assign rcache_line[7][54].status_reg.re    = reg2hw.status_1846.re;


  assign rcache_line[7][55].tag_reg.tag      = reg2hw.tag_1847.q;
  assign rcache_line[7][55].tag_reg.qe       = reg2hw.tag_1847.qe;
  assign rcache_line[7][55].tag_reg.re       = reg2hw.tag_1847.re;
  assign rcache_line[7][55].status_reg.status = reg2hw.status_1847.q;//status_reg_t'(reg2hw.status_1847.q);
  assign rcache_line[7][55].status_reg.qe    = reg2hw.status_1847.qe;
  assign rcache_line[7][55].status_reg.re    = reg2hw.status_1847.re;


  assign rcache_line[7][56].tag_reg.tag      = reg2hw.tag_1848.q;
  assign rcache_line[7][56].tag_reg.qe       = reg2hw.tag_1848.qe;
  assign rcache_line[7][56].tag_reg.re       = reg2hw.tag_1848.re;
  assign rcache_line[7][56].status_reg.status = reg2hw.status_1848.q;//status_reg_t'(reg2hw.status_1848.q);
  assign rcache_line[7][56].status_reg.qe    = reg2hw.status_1848.qe;
  assign rcache_line[7][56].status_reg.re    = reg2hw.status_1848.re;


  assign rcache_line[7][57].tag_reg.tag      = reg2hw.tag_1849.q;
  assign rcache_line[7][57].tag_reg.qe       = reg2hw.tag_1849.qe;
  assign rcache_line[7][57].tag_reg.re       = reg2hw.tag_1849.re;
  assign rcache_line[7][57].status_reg.status = reg2hw.status_1849.q;//status_reg_t'(reg2hw.status_1849.q);
  assign rcache_line[7][57].status_reg.qe    = reg2hw.status_1849.qe;
  assign rcache_line[7][57].status_reg.re    = reg2hw.status_1849.re;


  assign rcache_line[7][58].tag_reg.tag      = reg2hw.tag_1850.q;
  assign rcache_line[7][58].tag_reg.qe       = reg2hw.tag_1850.qe;
  assign rcache_line[7][58].tag_reg.re       = reg2hw.tag_1850.re;
  assign rcache_line[7][58].status_reg.status = reg2hw.status_1850.q;//status_reg_t'(reg2hw.status_1850.q);
  assign rcache_line[7][58].status_reg.qe    = reg2hw.status_1850.qe;
  assign rcache_line[7][58].status_reg.re    = reg2hw.status_1850.re;


  assign rcache_line[7][59].tag_reg.tag      = reg2hw.tag_1851.q;
  assign rcache_line[7][59].tag_reg.qe       = reg2hw.tag_1851.qe;
  assign rcache_line[7][59].tag_reg.re       = reg2hw.tag_1851.re;
  assign rcache_line[7][59].status_reg.status = reg2hw.status_1851.q;//status_reg_t'(reg2hw.status_1851.q);
  assign rcache_line[7][59].status_reg.qe    = reg2hw.status_1851.qe;
  assign rcache_line[7][59].status_reg.re    = reg2hw.status_1851.re;


  assign rcache_line[7][60].tag_reg.tag      = reg2hw.tag_1852.q;
  assign rcache_line[7][60].tag_reg.qe       = reg2hw.tag_1852.qe;
  assign rcache_line[7][60].tag_reg.re       = reg2hw.tag_1852.re;
  assign rcache_line[7][60].status_reg.status = reg2hw.status_1852.q;//status_reg_t'(reg2hw.status_1852.q);
  assign rcache_line[7][60].status_reg.qe    = reg2hw.status_1852.qe;
  assign rcache_line[7][60].status_reg.re    = reg2hw.status_1852.re;


  assign rcache_line[7][61].tag_reg.tag      = reg2hw.tag_1853.q;
  assign rcache_line[7][61].tag_reg.qe       = reg2hw.tag_1853.qe;
  assign rcache_line[7][61].tag_reg.re       = reg2hw.tag_1853.re;
  assign rcache_line[7][61].status_reg.status = reg2hw.status_1853.q;//status_reg_t'(reg2hw.status_1853.q);
  assign rcache_line[7][61].status_reg.qe    = reg2hw.status_1853.qe;
  assign rcache_line[7][61].status_reg.re    = reg2hw.status_1853.re;


  assign rcache_line[7][62].tag_reg.tag      = reg2hw.tag_1854.q;
  assign rcache_line[7][62].tag_reg.qe       = reg2hw.tag_1854.qe;
  assign rcache_line[7][62].tag_reg.re       = reg2hw.tag_1854.re;
  assign rcache_line[7][62].status_reg.status = reg2hw.status_1854.q;//status_reg_t'(reg2hw.status_1854.q);
  assign rcache_line[7][62].status_reg.qe    = reg2hw.status_1854.qe;
  assign rcache_line[7][62].status_reg.re    = reg2hw.status_1854.re;


  assign rcache_line[7][63].tag_reg.tag      = reg2hw.tag_1855.q;
  assign rcache_line[7][63].tag_reg.qe       = reg2hw.tag_1855.qe;
  assign rcache_line[7][63].tag_reg.re       = reg2hw.tag_1855.re;
  assign rcache_line[7][63].status_reg.status = reg2hw.status_1855.q;//status_reg_t'(reg2hw.status_1855.q);
  assign rcache_line[7][63].status_reg.qe    = reg2hw.status_1855.qe;
  assign rcache_line[7][63].status_reg.re    = reg2hw.status_1855.re;


  assign rcache_line[7][64].tag_reg.tag      = reg2hw.tag_1856.q;
  assign rcache_line[7][64].tag_reg.qe       = reg2hw.tag_1856.qe;
  assign rcache_line[7][64].tag_reg.re       = reg2hw.tag_1856.re;
  assign rcache_line[7][64].status_reg.status = reg2hw.status_1856.q;//status_reg_t'(reg2hw.status_1856.q);
  assign rcache_line[7][64].status_reg.qe    = reg2hw.status_1856.qe;
  assign rcache_line[7][64].status_reg.re    = reg2hw.status_1856.re;


  assign rcache_line[7][65].tag_reg.tag      = reg2hw.tag_1857.q;
  assign rcache_line[7][65].tag_reg.qe       = reg2hw.tag_1857.qe;
  assign rcache_line[7][65].tag_reg.re       = reg2hw.tag_1857.re;
  assign rcache_line[7][65].status_reg.status = reg2hw.status_1857.q;//status_reg_t'(reg2hw.status_1857.q);
  assign rcache_line[7][65].status_reg.qe    = reg2hw.status_1857.qe;
  assign rcache_line[7][65].status_reg.re    = reg2hw.status_1857.re;


  assign rcache_line[7][66].tag_reg.tag      = reg2hw.tag_1858.q;
  assign rcache_line[7][66].tag_reg.qe       = reg2hw.tag_1858.qe;
  assign rcache_line[7][66].tag_reg.re       = reg2hw.tag_1858.re;
  assign rcache_line[7][66].status_reg.status = reg2hw.status_1858.q;//status_reg_t'(reg2hw.status_1858.q);
  assign rcache_line[7][66].status_reg.qe    = reg2hw.status_1858.qe;
  assign rcache_line[7][66].status_reg.re    = reg2hw.status_1858.re;


  assign rcache_line[7][67].tag_reg.tag      = reg2hw.tag_1859.q;
  assign rcache_line[7][67].tag_reg.qe       = reg2hw.tag_1859.qe;
  assign rcache_line[7][67].tag_reg.re       = reg2hw.tag_1859.re;
  assign rcache_line[7][67].status_reg.status = reg2hw.status_1859.q;//status_reg_t'(reg2hw.status_1859.q);
  assign rcache_line[7][67].status_reg.qe    = reg2hw.status_1859.qe;
  assign rcache_line[7][67].status_reg.re    = reg2hw.status_1859.re;


  assign rcache_line[7][68].tag_reg.tag      = reg2hw.tag_1860.q;
  assign rcache_line[7][68].tag_reg.qe       = reg2hw.tag_1860.qe;
  assign rcache_line[7][68].tag_reg.re       = reg2hw.tag_1860.re;
  assign rcache_line[7][68].status_reg.status = reg2hw.status_1860.q;//status_reg_t'(reg2hw.status_1860.q);
  assign rcache_line[7][68].status_reg.qe    = reg2hw.status_1860.qe;
  assign rcache_line[7][68].status_reg.re    = reg2hw.status_1860.re;


  assign rcache_line[7][69].tag_reg.tag      = reg2hw.tag_1861.q;
  assign rcache_line[7][69].tag_reg.qe       = reg2hw.tag_1861.qe;
  assign rcache_line[7][69].tag_reg.re       = reg2hw.tag_1861.re;
  assign rcache_line[7][69].status_reg.status = reg2hw.status_1861.q;//status_reg_t'(reg2hw.status_1861.q);
  assign rcache_line[7][69].status_reg.qe    = reg2hw.status_1861.qe;
  assign rcache_line[7][69].status_reg.re    = reg2hw.status_1861.re;


  assign rcache_line[7][70].tag_reg.tag      = reg2hw.tag_1862.q;
  assign rcache_line[7][70].tag_reg.qe       = reg2hw.tag_1862.qe;
  assign rcache_line[7][70].tag_reg.re       = reg2hw.tag_1862.re;
  assign rcache_line[7][70].status_reg.status = reg2hw.status_1862.q;//status_reg_t'(reg2hw.status_1862.q);
  assign rcache_line[7][70].status_reg.qe    = reg2hw.status_1862.qe;
  assign rcache_line[7][70].status_reg.re    = reg2hw.status_1862.re;


  assign rcache_line[7][71].tag_reg.tag      = reg2hw.tag_1863.q;
  assign rcache_line[7][71].tag_reg.qe       = reg2hw.tag_1863.qe;
  assign rcache_line[7][71].tag_reg.re       = reg2hw.tag_1863.re;
  assign rcache_line[7][71].status_reg.status = reg2hw.status_1863.q;//status_reg_t'(reg2hw.status_1863.q);
  assign rcache_line[7][71].status_reg.qe    = reg2hw.status_1863.qe;
  assign rcache_line[7][71].status_reg.re    = reg2hw.status_1863.re;


  assign rcache_line[7][72].tag_reg.tag      = reg2hw.tag_1864.q;
  assign rcache_line[7][72].tag_reg.qe       = reg2hw.tag_1864.qe;
  assign rcache_line[7][72].tag_reg.re       = reg2hw.tag_1864.re;
  assign rcache_line[7][72].status_reg.status = reg2hw.status_1864.q;//status_reg_t'(reg2hw.status_1864.q);
  assign rcache_line[7][72].status_reg.qe    = reg2hw.status_1864.qe;
  assign rcache_line[7][72].status_reg.re    = reg2hw.status_1864.re;


  assign rcache_line[7][73].tag_reg.tag      = reg2hw.tag_1865.q;
  assign rcache_line[7][73].tag_reg.qe       = reg2hw.tag_1865.qe;
  assign rcache_line[7][73].tag_reg.re       = reg2hw.tag_1865.re;
  assign rcache_line[7][73].status_reg.status = reg2hw.status_1865.q;//status_reg_t'(reg2hw.status_1865.q);
  assign rcache_line[7][73].status_reg.qe    = reg2hw.status_1865.qe;
  assign rcache_line[7][73].status_reg.re    = reg2hw.status_1865.re;


  assign rcache_line[7][74].tag_reg.tag      = reg2hw.tag_1866.q;
  assign rcache_line[7][74].tag_reg.qe       = reg2hw.tag_1866.qe;
  assign rcache_line[7][74].tag_reg.re       = reg2hw.tag_1866.re;
  assign rcache_line[7][74].status_reg.status = reg2hw.status_1866.q;//status_reg_t'(reg2hw.status_1866.q);
  assign rcache_line[7][74].status_reg.qe    = reg2hw.status_1866.qe;
  assign rcache_line[7][74].status_reg.re    = reg2hw.status_1866.re;


  assign rcache_line[7][75].tag_reg.tag      = reg2hw.tag_1867.q;
  assign rcache_line[7][75].tag_reg.qe       = reg2hw.tag_1867.qe;
  assign rcache_line[7][75].tag_reg.re       = reg2hw.tag_1867.re;
  assign rcache_line[7][75].status_reg.status = reg2hw.status_1867.q;//status_reg_t'(reg2hw.status_1867.q);
  assign rcache_line[7][75].status_reg.qe    = reg2hw.status_1867.qe;
  assign rcache_line[7][75].status_reg.re    = reg2hw.status_1867.re;


  assign rcache_line[7][76].tag_reg.tag      = reg2hw.tag_1868.q;
  assign rcache_line[7][76].tag_reg.qe       = reg2hw.tag_1868.qe;
  assign rcache_line[7][76].tag_reg.re       = reg2hw.tag_1868.re;
  assign rcache_line[7][76].status_reg.status = reg2hw.status_1868.q;//status_reg_t'(reg2hw.status_1868.q);
  assign rcache_line[7][76].status_reg.qe    = reg2hw.status_1868.qe;
  assign rcache_line[7][76].status_reg.re    = reg2hw.status_1868.re;


  assign rcache_line[7][77].tag_reg.tag      = reg2hw.tag_1869.q;
  assign rcache_line[7][77].tag_reg.qe       = reg2hw.tag_1869.qe;
  assign rcache_line[7][77].tag_reg.re       = reg2hw.tag_1869.re;
  assign rcache_line[7][77].status_reg.status = reg2hw.status_1869.q;//status_reg_t'(reg2hw.status_1869.q);
  assign rcache_line[7][77].status_reg.qe    = reg2hw.status_1869.qe;
  assign rcache_line[7][77].status_reg.re    = reg2hw.status_1869.re;


  assign rcache_line[7][78].tag_reg.tag      = reg2hw.tag_1870.q;
  assign rcache_line[7][78].tag_reg.qe       = reg2hw.tag_1870.qe;
  assign rcache_line[7][78].tag_reg.re       = reg2hw.tag_1870.re;
  assign rcache_line[7][78].status_reg.status = reg2hw.status_1870.q;//status_reg_t'(reg2hw.status_1870.q);
  assign rcache_line[7][78].status_reg.qe    = reg2hw.status_1870.qe;
  assign rcache_line[7][78].status_reg.re    = reg2hw.status_1870.re;


  assign rcache_line[7][79].tag_reg.tag      = reg2hw.tag_1871.q;
  assign rcache_line[7][79].tag_reg.qe       = reg2hw.tag_1871.qe;
  assign rcache_line[7][79].tag_reg.re       = reg2hw.tag_1871.re;
  assign rcache_line[7][79].status_reg.status = reg2hw.status_1871.q;//status_reg_t'(reg2hw.status_1871.q);
  assign rcache_line[7][79].status_reg.qe    = reg2hw.status_1871.qe;
  assign rcache_line[7][79].status_reg.re    = reg2hw.status_1871.re;


  assign rcache_line[7][80].tag_reg.tag      = reg2hw.tag_1872.q;
  assign rcache_line[7][80].tag_reg.qe       = reg2hw.tag_1872.qe;
  assign rcache_line[7][80].tag_reg.re       = reg2hw.tag_1872.re;
  assign rcache_line[7][80].status_reg.status = reg2hw.status_1872.q;//status_reg_t'(reg2hw.status_1872.q);
  assign rcache_line[7][80].status_reg.qe    = reg2hw.status_1872.qe;
  assign rcache_line[7][80].status_reg.re    = reg2hw.status_1872.re;


  assign rcache_line[7][81].tag_reg.tag      = reg2hw.tag_1873.q;
  assign rcache_line[7][81].tag_reg.qe       = reg2hw.tag_1873.qe;
  assign rcache_line[7][81].tag_reg.re       = reg2hw.tag_1873.re;
  assign rcache_line[7][81].status_reg.status = reg2hw.status_1873.q;//status_reg_t'(reg2hw.status_1873.q);
  assign rcache_line[7][81].status_reg.qe    = reg2hw.status_1873.qe;
  assign rcache_line[7][81].status_reg.re    = reg2hw.status_1873.re;


  assign rcache_line[7][82].tag_reg.tag      = reg2hw.tag_1874.q;
  assign rcache_line[7][82].tag_reg.qe       = reg2hw.tag_1874.qe;
  assign rcache_line[7][82].tag_reg.re       = reg2hw.tag_1874.re;
  assign rcache_line[7][82].status_reg.status = reg2hw.status_1874.q;//status_reg_t'(reg2hw.status_1874.q);
  assign rcache_line[7][82].status_reg.qe    = reg2hw.status_1874.qe;
  assign rcache_line[7][82].status_reg.re    = reg2hw.status_1874.re;


  assign rcache_line[7][83].tag_reg.tag      = reg2hw.tag_1875.q;
  assign rcache_line[7][83].tag_reg.qe       = reg2hw.tag_1875.qe;
  assign rcache_line[7][83].tag_reg.re       = reg2hw.tag_1875.re;
  assign rcache_line[7][83].status_reg.status = reg2hw.status_1875.q;//status_reg_t'(reg2hw.status_1875.q);
  assign rcache_line[7][83].status_reg.qe    = reg2hw.status_1875.qe;
  assign rcache_line[7][83].status_reg.re    = reg2hw.status_1875.re;


  assign rcache_line[7][84].tag_reg.tag      = reg2hw.tag_1876.q;
  assign rcache_line[7][84].tag_reg.qe       = reg2hw.tag_1876.qe;
  assign rcache_line[7][84].tag_reg.re       = reg2hw.tag_1876.re;
  assign rcache_line[7][84].status_reg.status = reg2hw.status_1876.q;//status_reg_t'(reg2hw.status_1876.q);
  assign rcache_line[7][84].status_reg.qe    = reg2hw.status_1876.qe;
  assign rcache_line[7][84].status_reg.re    = reg2hw.status_1876.re;


  assign rcache_line[7][85].tag_reg.tag      = reg2hw.tag_1877.q;
  assign rcache_line[7][85].tag_reg.qe       = reg2hw.tag_1877.qe;
  assign rcache_line[7][85].tag_reg.re       = reg2hw.tag_1877.re;
  assign rcache_line[7][85].status_reg.status = reg2hw.status_1877.q;//status_reg_t'(reg2hw.status_1877.q);
  assign rcache_line[7][85].status_reg.qe    = reg2hw.status_1877.qe;
  assign rcache_line[7][85].status_reg.re    = reg2hw.status_1877.re;


  assign rcache_line[7][86].tag_reg.tag      = reg2hw.tag_1878.q;
  assign rcache_line[7][86].tag_reg.qe       = reg2hw.tag_1878.qe;
  assign rcache_line[7][86].tag_reg.re       = reg2hw.tag_1878.re;
  assign rcache_line[7][86].status_reg.status = reg2hw.status_1878.q;//status_reg_t'(reg2hw.status_1878.q);
  assign rcache_line[7][86].status_reg.qe    = reg2hw.status_1878.qe;
  assign rcache_line[7][86].status_reg.re    = reg2hw.status_1878.re;


  assign rcache_line[7][87].tag_reg.tag      = reg2hw.tag_1879.q;
  assign rcache_line[7][87].tag_reg.qe       = reg2hw.tag_1879.qe;
  assign rcache_line[7][87].tag_reg.re       = reg2hw.tag_1879.re;
  assign rcache_line[7][87].status_reg.status = reg2hw.status_1879.q;//status_reg_t'(reg2hw.status_1879.q);
  assign rcache_line[7][87].status_reg.qe    = reg2hw.status_1879.qe;
  assign rcache_line[7][87].status_reg.re    = reg2hw.status_1879.re;


  assign rcache_line[7][88].tag_reg.tag      = reg2hw.tag_1880.q;
  assign rcache_line[7][88].tag_reg.qe       = reg2hw.tag_1880.qe;
  assign rcache_line[7][88].tag_reg.re       = reg2hw.tag_1880.re;
  assign rcache_line[7][88].status_reg.status = reg2hw.status_1880.q;//status_reg_t'(reg2hw.status_1880.q);
  assign rcache_line[7][88].status_reg.qe    = reg2hw.status_1880.qe;
  assign rcache_line[7][88].status_reg.re    = reg2hw.status_1880.re;


  assign rcache_line[7][89].tag_reg.tag      = reg2hw.tag_1881.q;
  assign rcache_line[7][89].tag_reg.qe       = reg2hw.tag_1881.qe;
  assign rcache_line[7][89].tag_reg.re       = reg2hw.tag_1881.re;
  assign rcache_line[7][89].status_reg.status = reg2hw.status_1881.q;//status_reg_t'(reg2hw.status_1881.q);
  assign rcache_line[7][89].status_reg.qe    = reg2hw.status_1881.qe;
  assign rcache_line[7][89].status_reg.re    = reg2hw.status_1881.re;


  assign rcache_line[7][90].tag_reg.tag      = reg2hw.tag_1882.q;
  assign rcache_line[7][90].tag_reg.qe       = reg2hw.tag_1882.qe;
  assign rcache_line[7][90].tag_reg.re       = reg2hw.tag_1882.re;
  assign rcache_line[7][90].status_reg.status = reg2hw.status_1882.q;//status_reg_t'(reg2hw.status_1882.q);
  assign rcache_line[7][90].status_reg.qe    = reg2hw.status_1882.qe;
  assign rcache_line[7][90].status_reg.re    = reg2hw.status_1882.re;


  assign rcache_line[7][91].tag_reg.tag      = reg2hw.tag_1883.q;
  assign rcache_line[7][91].tag_reg.qe       = reg2hw.tag_1883.qe;
  assign rcache_line[7][91].tag_reg.re       = reg2hw.tag_1883.re;
  assign rcache_line[7][91].status_reg.status = reg2hw.status_1883.q;//status_reg_t'(reg2hw.status_1883.q);
  assign rcache_line[7][91].status_reg.qe    = reg2hw.status_1883.qe;
  assign rcache_line[7][91].status_reg.re    = reg2hw.status_1883.re;


  assign rcache_line[7][92].tag_reg.tag      = reg2hw.tag_1884.q;
  assign rcache_line[7][92].tag_reg.qe       = reg2hw.tag_1884.qe;
  assign rcache_line[7][92].tag_reg.re       = reg2hw.tag_1884.re;
  assign rcache_line[7][92].status_reg.status = reg2hw.status_1884.q;//status_reg_t'(reg2hw.status_1884.q);
  assign rcache_line[7][92].status_reg.qe    = reg2hw.status_1884.qe;
  assign rcache_line[7][92].status_reg.re    = reg2hw.status_1884.re;


  assign rcache_line[7][93].tag_reg.tag      = reg2hw.tag_1885.q;
  assign rcache_line[7][93].tag_reg.qe       = reg2hw.tag_1885.qe;
  assign rcache_line[7][93].tag_reg.re       = reg2hw.tag_1885.re;
  assign rcache_line[7][93].status_reg.status = reg2hw.status_1885.q;//status_reg_t'(reg2hw.status_1885.q);
  assign rcache_line[7][93].status_reg.qe    = reg2hw.status_1885.qe;
  assign rcache_line[7][93].status_reg.re    = reg2hw.status_1885.re;


  assign rcache_line[7][94].tag_reg.tag      = reg2hw.tag_1886.q;
  assign rcache_line[7][94].tag_reg.qe       = reg2hw.tag_1886.qe;
  assign rcache_line[7][94].tag_reg.re       = reg2hw.tag_1886.re;
  assign rcache_line[7][94].status_reg.status = reg2hw.status_1886.q;//status_reg_t'(reg2hw.status_1886.q);
  assign rcache_line[7][94].status_reg.qe    = reg2hw.status_1886.qe;
  assign rcache_line[7][94].status_reg.re    = reg2hw.status_1886.re;


  assign rcache_line[7][95].tag_reg.tag      = reg2hw.tag_1887.q;
  assign rcache_line[7][95].tag_reg.qe       = reg2hw.tag_1887.qe;
  assign rcache_line[7][95].tag_reg.re       = reg2hw.tag_1887.re;
  assign rcache_line[7][95].status_reg.status = reg2hw.status_1887.q;//status_reg_t'(reg2hw.status_1887.q);
  assign rcache_line[7][95].status_reg.qe    = reg2hw.status_1887.qe;
  assign rcache_line[7][95].status_reg.re    = reg2hw.status_1887.re;


  assign rcache_line[7][96].tag_reg.tag      = reg2hw.tag_1888.q;
  assign rcache_line[7][96].tag_reg.qe       = reg2hw.tag_1888.qe;
  assign rcache_line[7][96].tag_reg.re       = reg2hw.tag_1888.re;
  assign rcache_line[7][96].status_reg.status = reg2hw.status_1888.q;//status_reg_t'(reg2hw.status_1888.q);
  assign rcache_line[7][96].status_reg.qe    = reg2hw.status_1888.qe;
  assign rcache_line[7][96].status_reg.re    = reg2hw.status_1888.re;


  assign rcache_line[7][97].tag_reg.tag      = reg2hw.tag_1889.q;
  assign rcache_line[7][97].tag_reg.qe       = reg2hw.tag_1889.qe;
  assign rcache_line[7][97].tag_reg.re       = reg2hw.tag_1889.re;
  assign rcache_line[7][97].status_reg.status = reg2hw.status_1889.q;//status_reg_t'(reg2hw.status_1889.q);
  assign rcache_line[7][97].status_reg.qe    = reg2hw.status_1889.qe;
  assign rcache_line[7][97].status_reg.re    = reg2hw.status_1889.re;


  assign rcache_line[7][98].tag_reg.tag      = reg2hw.tag_1890.q;
  assign rcache_line[7][98].tag_reg.qe       = reg2hw.tag_1890.qe;
  assign rcache_line[7][98].tag_reg.re       = reg2hw.tag_1890.re;
  assign rcache_line[7][98].status_reg.status = reg2hw.status_1890.q;//status_reg_t'(reg2hw.status_1890.q);
  assign rcache_line[7][98].status_reg.qe    = reg2hw.status_1890.qe;
  assign rcache_line[7][98].status_reg.re    = reg2hw.status_1890.re;


  assign rcache_line[7][99].tag_reg.tag      = reg2hw.tag_1891.q;
  assign rcache_line[7][99].tag_reg.qe       = reg2hw.tag_1891.qe;
  assign rcache_line[7][99].tag_reg.re       = reg2hw.tag_1891.re;
  assign rcache_line[7][99].status_reg.status = reg2hw.status_1891.q;//status_reg_t'(reg2hw.status_1891.q);
  assign rcache_line[7][99].status_reg.qe    = reg2hw.status_1891.qe;
  assign rcache_line[7][99].status_reg.re    = reg2hw.status_1891.re;


  assign rcache_line[7][100].tag_reg.tag      = reg2hw.tag_1892.q;
  assign rcache_line[7][100].tag_reg.qe       = reg2hw.tag_1892.qe;
  assign rcache_line[7][100].tag_reg.re       = reg2hw.tag_1892.re;
  assign rcache_line[7][100].status_reg.status = reg2hw.status_1892.q;//status_reg_t'(reg2hw.status_1892.q);
  assign rcache_line[7][100].status_reg.qe    = reg2hw.status_1892.qe;
  assign rcache_line[7][100].status_reg.re    = reg2hw.status_1892.re;


  assign rcache_line[7][101].tag_reg.tag      = reg2hw.tag_1893.q;
  assign rcache_line[7][101].tag_reg.qe       = reg2hw.tag_1893.qe;
  assign rcache_line[7][101].tag_reg.re       = reg2hw.tag_1893.re;
  assign rcache_line[7][101].status_reg.status = reg2hw.status_1893.q;//status_reg_t'(reg2hw.status_1893.q);
  assign rcache_line[7][101].status_reg.qe    = reg2hw.status_1893.qe;
  assign rcache_line[7][101].status_reg.re    = reg2hw.status_1893.re;


  assign rcache_line[7][102].tag_reg.tag      = reg2hw.tag_1894.q;
  assign rcache_line[7][102].tag_reg.qe       = reg2hw.tag_1894.qe;
  assign rcache_line[7][102].tag_reg.re       = reg2hw.tag_1894.re;
  assign rcache_line[7][102].status_reg.status = reg2hw.status_1894.q;//status_reg_t'(reg2hw.status_1894.q);
  assign rcache_line[7][102].status_reg.qe    = reg2hw.status_1894.qe;
  assign rcache_line[7][102].status_reg.re    = reg2hw.status_1894.re;


  assign rcache_line[7][103].tag_reg.tag      = reg2hw.tag_1895.q;
  assign rcache_line[7][103].tag_reg.qe       = reg2hw.tag_1895.qe;
  assign rcache_line[7][103].tag_reg.re       = reg2hw.tag_1895.re;
  assign rcache_line[7][103].status_reg.status = reg2hw.status_1895.q;//status_reg_t'(reg2hw.status_1895.q);
  assign rcache_line[7][103].status_reg.qe    = reg2hw.status_1895.qe;
  assign rcache_line[7][103].status_reg.re    = reg2hw.status_1895.re;


  assign rcache_line[7][104].tag_reg.tag      = reg2hw.tag_1896.q;
  assign rcache_line[7][104].tag_reg.qe       = reg2hw.tag_1896.qe;
  assign rcache_line[7][104].tag_reg.re       = reg2hw.tag_1896.re;
  assign rcache_line[7][104].status_reg.status = reg2hw.status_1896.q;//status_reg_t'(reg2hw.status_1896.q);
  assign rcache_line[7][104].status_reg.qe    = reg2hw.status_1896.qe;
  assign rcache_line[7][104].status_reg.re    = reg2hw.status_1896.re;


  assign rcache_line[7][105].tag_reg.tag      = reg2hw.tag_1897.q;
  assign rcache_line[7][105].tag_reg.qe       = reg2hw.tag_1897.qe;
  assign rcache_line[7][105].tag_reg.re       = reg2hw.tag_1897.re;
  assign rcache_line[7][105].status_reg.status = reg2hw.status_1897.q;//status_reg_t'(reg2hw.status_1897.q);
  assign rcache_line[7][105].status_reg.qe    = reg2hw.status_1897.qe;
  assign rcache_line[7][105].status_reg.re    = reg2hw.status_1897.re;


  assign rcache_line[7][106].tag_reg.tag      = reg2hw.tag_1898.q;
  assign rcache_line[7][106].tag_reg.qe       = reg2hw.tag_1898.qe;
  assign rcache_line[7][106].tag_reg.re       = reg2hw.tag_1898.re;
  assign rcache_line[7][106].status_reg.status = reg2hw.status_1898.q;//status_reg_t'(reg2hw.status_1898.q);
  assign rcache_line[7][106].status_reg.qe    = reg2hw.status_1898.qe;
  assign rcache_line[7][106].status_reg.re    = reg2hw.status_1898.re;


  assign rcache_line[7][107].tag_reg.tag      = reg2hw.tag_1899.q;
  assign rcache_line[7][107].tag_reg.qe       = reg2hw.tag_1899.qe;
  assign rcache_line[7][107].tag_reg.re       = reg2hw.tag_1899.re;
  assign rcache_line[7][107].status_reg.status = reg2hw.status_1899.q;//status_reg_t'(reg2hw.status_1899.q);
  assign rcache_line[7][107].status_reg.qe    = reg2hw.status_1899.qe;
  assign rcache_line[7][107].status_reg.re    = reg2hw.status_1899.re;


  assign rcache_line[7][108].tag_reg.tag      = reg2hw.tag_1900.q;
  assign rcache_line[7][108].tag_reg.qe       = reg2hw.tag_1900.qe;
  assign rcache_line[7][108].tag_reg.re       = reg2hw.tag_1900.re;
  assign rcache_line[7][108].status_reg.status = reg2hw.status_1900.q;//status_reg_t'(reg2hw.status_1900.q);
  assign rcache_line[7][108].status_reg.qe    = reg2hw.status_1900.qe;
  assign rcache_line[7][108].status_reg.re    = reg2hw.status_1900.re;


  assign rcache_line[7][109].tag_reg.tag      = reg2hw.tag_1901.q;
  assign rcache_line[7][109].tag_reg.qe       = reg2hw.tag_1901.qe;
  assign rcache_line[7][109].tag_reg.re       = reg2hw.tag_1901.re;
  assign rcache_line[7][109].status_reg.status = reg2hw.status_1901.q;//status_reg_t'(reg2hw.status_1901.q);
  assign rcache_line[7][109].status_reg.qe    = reg2hw.status_1901.qe;
  assign rcache_line[7][109].status_reg.re    = reg2hw.status_1901.re;


  assign rcache_line[7][110].tag_reg.tag      = reg2hw.tag_1902.q;
  assign rcache_line[7][110].tag_reg.qe       = reg2hw.tag_1902.qe;
  assign rcache_line[7][110].tag_reg.re       = reg2hw.tag_1902.re;
  assign rcache_line[7][110].status_reg.status = reg2hw.status_1902.q;//status_reg_t'(reg2hw.status_1902.q);
  assign rcache_line[7][110].status_reg.qe    = reg2hw.status_1902.qe;
  assign rcache_line[7][110].status_reg.re    = reg2hw.status_1902.re;


  assign rcache_line[7][111].tag_reg.tag      = reg2hw.tag_1903.q;
  assign rcache_line[7][111].tag_reg.qe       = reg2hw.tag_1903.qe;
  assign rcache_line[7][111].tag_reg.re       = reg2hw.tag_1903.re;
  assign rcache_line[7][111].status_reg.status = reg2hw.status_1903.q;//status_reg_t'(reg2hw.status_1903.q);
  assign rcache_line[7][111].status_reg.qe    = reg2hw.status_1903.qe;
  assign rcache_line[7][111].status_reg.re    = reg2hw.status_1903.re;


  assign rcache_line[7][112].tag_reg.tag      = reg2hw.tag_1904.q;
  assign rcache_line[7][112].tag_reg.qe       = reg2hw.tag_1904.qe;
  assign rcache_line[7][112].tag_reg.re       = reg2hw.tag_1904.re;
  assign rcache_line[7][112].status_reg.status = reg2hw.status_1904.q;//status_reg_t'(reg2hw.status_1904.q);
  assign rcache_line[7][112].status_reg.qe    = reg2hw.status_1904.qe;
  assign rcache_line[7][112].status_reg.re    = reg2hw.status_1904.re;


  assign rcache_line[7][113].tag_reg.tag      = reg2hw.tag_1905.q;
  assign rcache_line[7][113].tag_reg.qe       = reg2hw.tag_1905.qe;
  assign rcache_line[7][113].tag_reg.re       = reg2hw.tag_1905.re;
  assign rcache_line[7][113].status_reg.status = reg2hw.status_1905.q;//status_reg_t'(reg2hw.status_1905.q);
  assign rcache_line[7][113].status_reg.qe    = reg2hw.status_1905.qe;
  assign rcache_line[7][113].status_reg.re    = reg2hw.status_1905.re;


  assign rcache_line[7][114].tag_reg.tag      = reg2hw.tag_1906.q;
  assign rcache_line[7][114].tag_reg.qe       = reg2hw.tag_1906.qe;
  assign rcache_line[7][114].tag_reg.re       = reg2hw.tag_1906.re;
  assign rcache_line[7][114].status_reg.status = reg2hw.status_1906.q;//status_reg_t'(reg2hw.status_1906.q);
  assign rcache_line[7][114].status_reg.qe    = reg2hw.status_1906.qe;
  assign rcache_line[7][114].status_reg.re    = reg2hw.status_1906.re;


  assign rcache_line[7][115].tag_reg.tag      = reg2hw.tag_1907.q;
  assign rcache_line[7][115].tag_reg.qe       = reg2hw.tag_1907.qe;
  assign rcache_line[7][115].tag_reg.re       = reg2hw.tag_1907.re;
  assign rcache_line[7][115].status_reg.status = reg2hw.status_1907.q;//status_reg_t'(reg2hw.status_1907.q);
  assign rcache_line[7][115].status_reg.qe    = reg2hw.status_1907.qe;
  assign rcache_line[7][115].status_reg.re    = reg2hw.status_1907.re;


  assign rcache_line[7][116].tag_reg.tag      = reg2hw.tag_1908.q;
  assign rcache_line[7][116].tag_reg.qe       = reg2hw.tag_1908.qe;
  assign rcache_line[7][116].tag_reg.re       = reg2hw.tag_1908.re;
  assign rcache_line[7][116].status_reg.status = reg2hw.status_1908.q;//status_reg_t'(reg2hw.status_1908.q);
  assign rcache_line[7][116].status_reg.qe    = reg2hw.status_1908.qe;
  assign rcache_line[7][116].status_reg.re    = reg2hw.status_1908.re;


  assign rcache_line[7][117].tag_reg.tag      = reg2hw.tag_1909.q;
  assign rcache_line[7][117].tag_reg.qe       = reg2hw.tag_1909.qe;
  assign rcache_line[7][117].tag_reg.re       = reg2hw.tag_1909.re;
  assign rcache_line[7][117].status_reg.status = reg2hw.status_1909.q;//status_reg_t'(reg2hw.status_1909.q);
  assign rcache_line[7][117].status_reg.qe    = reg2hw.status_1909.qe;
  assign rcache_line[7][117].status_reg.re    = reg2hw.status_1909.re;


  assign rcache_line[7][118].tag_reg.tag      = reg2hw.tag_1910.q;
  assign rcache_line[7][118].tag_reg.qe       = reg2hw.tag_1910.qe;
  assign rcache_line[7][118].tag_reg.re       = reg2hw.tag_1910.re;
  assign rcache_line[7][118].status_reg.status = reg2hw.status_1910.q;//status_reg_t'(reg2hw.status_1910.q);
  assign rcache_line[7][118].status_reg.qe    = reg2hw.status_1910.qe;
  assign rcache_line[7][118].status_reg.re    = reg2hw.status_1910.re;


  assign rcache_line[7][119].tag_reg.tag      = reg2hw.tag_1911.q;
  assign rcache_line[7][119].tag_reg.qe       = reg2hw.tag_1911.qe;
  assign rcache_line[7][119].tag_reg.re       = reg2hw.tag_1911.re;
  assign rcache_line[7][119].status_reg.status = reg2hw.status_1911.q;//status_reg_t'(reg2hw.status_1911.q);
  assign rcache_line[7][119].status_reg.qe    = reg2hw.status_1911.qe;
  assign rcache_line[7][119].status_reg.re    = reg2hw.status_1911.re;


  assign rcache_line[7][120].tag_reg.tag      = reg2hw.tag_1912.q;
  assign rcache_line[7][120].tag_reg.qe       = reg2hw.tag_1912.qe;
  assign rcache_line[7][120].tag_reg.re       = reg2hw.tag_1912.re;
  assign rcache_line[7][120].status_reg.status = reg2hw.status_1912.q;//status_reg_t'(reg2hw.status_1912.q);
  assign rcache_line[7][120].status_reg.qe    = reg2hw.status_1912.qe;
  assign rcache_line[7][120].status_reg.re    = reg2hw.status_1912.re;


  assign rcache_line[7][121].tag_reg.tag      = reg2hw.tag_1913.q;
  assign rcache_line[7][121].tag_reg.qe       = reg2hw.tag_1913.qe;
  assign rcache_line[7][121].tag_reg.re       = reg2hw.tag_1913.re;
  assign rcache_line[7][121].status_reg.status = reg2hw.status_1913.q;//status_reg_t'(reg2hw.status_1913.q);
  assign rcache_line[7][121].status_reg.qe    = reg2hw.status_1913.qe;
  assign rcache_line[7][121].status_reg.re    = reg2hw.status_1913.re;


  assign rcache_line[7][122].tag_reg.tag      = reg2hw.tag_1914.q;
  assign rcache_line[7][122].tag_reg.qe       = reg2hw.tag_1914.qe;
  assign rcache_line[7][122].tag_reg.re       = reg2hw.tag_1914.re;
  assign rcache_line[7][122].status_reg.status = reg2hw.status_1914.q;//status_reg_t'(reg2hw.status_1914.q);
  assign rcache_line[7][122].status_reg.qe    = reg2hw.status_1914.qe;
  assign rcache_line[7][122].status_reg.re    = reg2hw.status_1914.re;


  assign rcache_line[7][123].tag_reg.tag      = reg2hw.tag_1915.q;
  assign rcache_line[7][123].tag_reg.qe       = reg2hw.tag_1915.qe;
  assign rcache_line[7][123].tag_reg.re       = reg2hw.tag_1915.re;
  assign rcache_line[7][123].status_reg.status = reg2hw.status_1915.q;//status_reg_t'(reg2hw.status_1915.q);
  assign rcache_line[7][123].status_reg.qe    = reg2hw.status_1915.qe;
  assign rcache_line[7][123].status_reg.re    = reg2hw.status_1915.re;


  assign rcache_line[7][124].tag_reg.tag      = reg2hw.tag_1916.q;
  assign rcache_line[7][124].tag_reg.qe       = reg2hw.tag_1916.qe;
  assign rcache_line[7][124].tag_reg.re       = reg2hw.tag_1916.re;
  assign rcache_line[7][124].status_reg.status = reg2hw.status_1916.q;//status_reg_t'(reg2hw.status_1916.q);
  assign rcache_line[7][124].status_reg.qe    = reg2hw.status_1916.qe;
  assign rcache_line[7][124].status_reg.re    = reg2hw.status_1916.re;


  assign rcache_line[7][125].tag_reg.tag      = reg2hw.tag_1917.q;
  assign rcache_line[7][125].tag_reg.qe       = reg2hw.tag_1917.qe;
  assign rcache_line[7][125].tag_reg.re       = reg2hw.tag_1917.re;
  assign rcache_line[7][125].status_reg.status = reg2hw.status_1917.q;//status_reg_t'(reg2hw.status_1917.q);
  assign rcache_line[7][125].status_reg.qe    = reg2hw.status_1917.qe;
  assign rcache_line[7][125].status_reg.re    = reg2hw.status_1917.re;


  assign rcache_line[7][126].tag_reg.tag      = reg2hw.tag_1918.q;
  assign rcache_line[7][126].tag_reg.qe       = reg2hw.tag_1918.qe;
  assign rcache_line[7][126].tag_reg.re       = reg2hw.tag_1918.re;
  assign rcache_line[7][126].status_reg.status = reg2hw.status_1918.q;//status_reg_t'(reg2hw.status_1918.q);
  assign rcache_line[7][126].status_reg.qe    = reg2hw.status_1918.qe;
  assign rcache_line[7][126].status_reg.re    = reg2hw.status_1918.re;


  assign rcache_line[7][127].tag_reg.tag      = reg2hw.tag_1919.q;
  assign rcache_line[7][127].tag_reg.qe       = reg2hw.tag_1919.qe;
  assign rcache_line[7][127].tag_reg.re       = reg2hw.tag_1919.re;
  assign rcache_line[7][127].status_reg.status = reg2hw.status_1919.q;//status_reg_t'(reg2hw.status_1919.q);
  assign rcache_line[7][127].status_reg.qe    = reg2hw.status_1919.qe;
  assign rcache_line[7][127].status_reg.re    = reg2hw.status_1919.re;


  assign rcache_line[7][128].tag_reg.tag      = reg2hw.tag_1920.q;
  assign rcache_line[7][128].tag_reg.qe       = reg2hw.tag_1920.qe;
  assign rcache_line[7][128].tag_reg.re       = reg2hw.tag_1920.re;
  assign rcache_line[7][128].status_reg.status = reg2hw.status_1920.q;//status_reg_t'(reg2hw.status_1920.q);
  assign rcache_line[7][128].status_reg.qe    = reg2hw.status_1920.qe;
  assign rcache_line[7][128].status_reg.re    = reg2hw.status_1920.re;


  assign rcache_line[7][129].tag_reg.tag      = reg2hw.tag_1921.q;
  assign rcache_line[7][129].tag_reg.qe       = reg2hw.tag_1921.qe;
  assign rcache_line[7][129].tag_reg.re       = reg2hw.tag_1921.re;
  assign rcache_line[7][129].status_reg.status = reg2hw.status_1921.q;//status_reg_t'(reg2hw.status_1921.q);
  assign rcache_line[7][129].status_reg.qe    = reg2hw.status_1921.qe;
  assign rcache_line[7][129].status_reg.re    = reg2hw.status_1921.re;


  assign rcache_line[7][130].tag_reg.tag      = reg2hw.tag_1922.q;
  assign rcache_line[7][130].tag_reg.qe       = reg2hw.tag_1922.qe;
  assign rcache_line[7][130].tag_reg.re       = reg2hw.tag_1922.re;
  assign rcache_line[7][130].status_reg.status = reg2hw.status_1922.q;//status_reg_t'(reg2hw.status_1922.q);
  assign rcache_line[7][130].status_reg.qe    = reg2hw.status_1922.qe;
  assign rcache_line[7][130].status_reg.re    = reg2hw.status_1922.re;


  assign rcache_line[7][131].tag_reg.tag      = reg2hw.tag_1923.q;
  assign rcache_line[7][131].tag_reg.qe       = reg2hw.tag_1923.qe;
  assign rcache_line[7][131].tag_reg.re       = reg2hw.tag_1923.re;
  assign rcache_line[7][131].status_reg.status = reg2hw.status_1923.q;//status_reg_t'(reg2hw.status_1923.q);
  assign rcache_line[7][131].status_reg.qe    = reg2hw.status_1923.qe;
  assign rcache_line[7][131].status_reg.re    = reg2hw.status_1923.re;


  assign rcache_line[7][132].tag_reg.tag      = reg2hw.tag_1924.q;
  assign rcache_line[7][132].tag_reg.qe       = reg2hw.tag_1924.qe;
  assign rcache_line[7][132].tag_reg.re       = reg2hw.tag_1924.re;
  assign rcache_line[7][132].status_reg.status = reg2hw.status_1924.q;//status_reg_t'(reg2hw.status_1924.q);
  assign rcache_line[7][132].status_reg.qe    = reg2hw.status_1924.qe;
  assign rcache_line[7][132].status_reg.re    = reg2hw.status_1924.re;


  assign rcache_line[7][133].tag_reg.tag      = reg2hw.tag_1925.q;
  assign rcache_line[7][133].tag_reg.qe       = reg2hw.tag_1925.qe;
  assign rcache_line[7][133].tag_reg.re       = reg2hw.tag_1925.re;
  assign rcache_line[7][133].status_reg.status = reg2hw.status_1925.q;//status_reg_t'(reg2hw.status_1925.q);
  assign rcache_line[7][133].status_reg.qe    = reg2hw.status_1925.qe;
  assign rcache_line[7][133].status_reg.re    = reg2hw.status_1925.re;


  assign rcache_line[7][134].tag_reg.tag      = reg2hw.tag_1926.q;
  assign rcache_line[7][134].tag_reg.qe       = reg2hw.tag_1926.qe;
  assign rcache_line[7][134].tag_reg.re       = reg2hw.tag_1926.re;
  assign rcache_line[7][134].status_reg.status = reg2hw.status_1926.q;//status_reg_t'(reg2hw.status_1926.q);
  assign rcache_line[7][134].status_reg.qe    = reg2hw.status_1926.qe;
  assign rcache_line[7][134].status_reg.re    = reg2hw.status_1926.re;


  assign rcache_line[7][135].tag_reg.tag      = reg2hw.tag_1927.q;
  assign rcache_line[7][135].tag_reg.qe       = reg2hw.tag_1927.qe;
  assign rcache_line[7][135].tag_reg.re       = reg2hw.tag_1927.re;
  assign rcache_line[7][135].status_reg.status = reg2hw.status_1927.q;//status_reg_t'(reg2hw.status_1927.q);
  assign rcache_line[7][135].status_reg.qe    = reg2hw.status_1927.qe;
  assign rcache_line[7][135].status_reg.re    = reg2hw.status_1927.re;


  assign rcache_line[7][136].tag_reg.tag      = reg2hw.tag_1928.q;
  assign rcache_line[7][136].tag_reg.qe       = reg2hw.tag_1928.qe;
  assign rcache_line[7][136].tag_reg.re       = reg2hw.tag_1928.re;
  assign rcache_line[7][136].status_reg.status = reg2hw.status_1928.q;//status_reg_t'(reg2hw.status_1928.q);
  assign rcache_line[7][136].status_reg.qe    = reg2hw.status_1928.qe;
  assign rcache_line[7][136].status_reg.re    = reg2hw.status_1928.re;


  assign rcache_line[7][137].tag_reg.tag      = reg2hw.tag_1929.q;
  assign rcache_line[7][137].tag_reg.qe       = reg2hw.tag_1929.qe;
  assign rcache_line[7][137].tag_reg.re       = reg2hw.tag_1929.re;
  assign rcache_line[7][137].status_reg.status = reg2hw.status_1929.q;//status_reg_t'(reg2hw.status_1929.q);
  assign rcache_line[7][137].status_reg.qe    = reg2hw.status_1929.qe;
  assign rcache_line[7][137].status_reg.re    = reg2hw.status_1929.re;


  assign rcache_line[7][138].tag_reg.tag      = reg2hw.tag_1930.q;
  assign rcache_line[7][138].tag_reg.qe       = reg2hw.tag_1930.qe;
  assign rcache_line[7][138].tag_reg.re       = reg2hw.tag_1930.re;
  assign rcache_line[7][138].status_reg.status = reg2hw.status_1930.q;//status_reg_t'(reg2hw.status_1930.q);
  assign rcache_line[7][138].status_reg.qe    = reg2hw.status_1930.qe;
  assign rcache_line[7][138].status_reg.re    = reg2hw.status_1930.re;


  assign rcache_line[7][139].tag_reg.tag      = reg2hw.tag_1931.q;
  assign rcache_line[7][139].tag_reg.qe       = reg2hw.tag_1931.qe;
  assign rcache_line[7][139].tag_reg.re       = reg2hw.tag_1931.re;
  assign rcache_line[7][139].status_reg.status = reg2hw.status_1931.q;//status_reg_t'(reg2hw.status_1931.q);
  assign rcache_line[7][139].status_reg.qe    = reg2hw.status_1931.qe;
  assign rcache_line[7][139].status_reg.re    = reg2hw.status_1931.re;


  assign rcache_line[7][140].tag_reg.tag      = reg2hw.tag_1932.q;
  assign rcache_line[7][140].tag_reg.qe       = reg2hw.tag_1932.qe;
  assign rcache_line[7][140].tag_reg.re       = reg2hw.tag_1932.re;
  assign rcache_line[7][140].status_reg.status = reg2hw.status_1932.q;//status_reg_t'(reg2hw.status_1932.q);
  assign rcache_line[7][140].status_reg.qe    = reg2hw.status_1932.qe;
  assign rcache_line[7][140].status_reg.re    = reg2hw.status_1932.re;


  assign rcache_line[7][141].tag_reg.tag      = reg2hw.tag_1933.q;
  assign rcache_line[7][141].tag_reg.qe       = reg2hw.tag_1933.qe;
  assign rcache_line[7][141].tag_reg.re       = reg2hw.tag_1933.re;
  assign rcache_line[7][141].status_reg.status = reg2hw.status_1933.q;//status_reg_t'(reg2hw.status_1933.q);
  assign rcache_line[7][141].status_reg.qe    = reg2hw.status_1933.qe;
  assign rcache_line[7][141].status_reg.re    = reg2hw.status_1933.re;


  assign rcache_line[7][142].tag_reg.tag      = reg2hw.tag_1934.q;
  assign rcache_line[7][142].tag_reg.qe       = reg2hw.tag_1934.qe;
  assign rcache_line[7][142].tag_reg.re       = reg2hw.tag_1934.re;
  assign rcache_line[7][142].status_reg.status = reg2hw.status_1934.q;//status_reg_t'(reg2hw.status_1934.q);
  assign rcache_line[7][142].status_reg.qe    = reg2hw.status_1934.qe;
  assign rcache_line[7][142].status_reg.re    = reg2hw.status_1934.re;


  assign rcache_line[7][143].tag_reg.tag      = reg2hw.tag_1935.q;
  assign rcache_line[7][143].tag_reg.qe       = reg2hw.tag_1935.qe;
  assign rcache_line[7][143].tag_reg.re       = reg2hw.tag_1935.re;
  assign rcache_line[7][143].status_reg.status = reg2hw.status_1935.q;//status_reg_t'(reg2hw.status_1935.q);
  assign rcache_line[7][143].status_reg.qe    = reg2hw.status_1935.qe;
  assign rcache_line[7][143].status_reg.re    = reg2hw.status_1935.re;


  assign rcache_line[7][144].tag_reg.tag      = reg2hw.tag_1936.q;
  assign rcache_line[7][144].tag_reg.qe       = reg2hw.tag_1936.qe;
  assign rcache_line[7][144].tag_reg.re       = reg2hw.tag_1936.re;
  assign rcache_line[7][144].status_reg.status = reg2hw.status_1936.q;//status_reg_t'(reg2hw.status_1936.q);
  assign rcache_line[7][144].status_reg.qe    = reg2hw.status_1936.qe;
  assign rcache_line[7][144].status_reg.re    = reg2hw.status_1936.re;


  assign rcache_line[7][145].tag_reg.tag      = reg2hw.tag_1937.q;
  assign rcache_line[7][145].tag_reg.qe       = reg2hw.tag_1937.qe;
  assign rcache_line[7][145].tag_reg.re       = reg2hw.tag_1937.re;
  assign rcache_line[7][145].status_reg.status = reg2hw.status_1937.q;//status_reg_t'(reg2hw.status_1937.q);
  assign rcache_line[7][145].status_reg.qe    = reg2hw.status_1937.qe;
  assign rcache_line[7][145].status_reg.re    = reg2hw.status_1937.re;


  assign rcache_line[7][146].tag_reg.tag      = reg2hw.tag_1938.q;
  assign rcache_line[7][146].tag_reg.qe       = reg2hw.tag_1938.qe;
  assign rcache_line[7][146].tag_reg.re       = reg2hw.tag_1938.re;
  assign rcache_line[7][146].status_reg.status = reg2hw.status_1938.q;//status_reg_t'(reg2hw.status_1938.q);
  assign rcache_line[7][146].status_reg.qe    = reg2hw.status_1938.qe;
  assign rcache_line[7][146].status_reg.re    = reg2hw.status_1938.re;


  assign rcache_line[7][147].tag_reg.tag      = reg2hw.tag_1939.q;
  assign rcache_line[7][147].tag_reg.qe       = reg2hw.tag_1939.qe;
  assign rcache_line[7][147].tag_reg.re       = reg2hw.tag_1939.re;
  assign rcache_line[7][147].status_reg.status = reg2hw.status_1939.q;//status_reg_t'(reg2hw.status_1939.q);
  assign rcache_line[7][147].status_reg.qe    = reg2hw.status_1939.qe;
  assign rcache_line[7][147].status_reg.re    = reg2hw.status_1939.re;


  assign rcache_line[7][148].tag_reg.tag      = reg2hw.tag_1940.q;
  assign rcache_line[7][148].tag_reg.qe       = reg2hw.tag_1940.qe;
  assign rcache_line[7][148].tag_reg.re       = reg2hw.tag_1940.re;
  assign rcache_line[7][148].status_reg.status = reg2hw.status_1940.q;//status_reg_t'(reg2hw.status_1940.q);
  assign rcache_line[7][148].status_reg.qe    = reg2hw.status_1940.qe;
  assign rcache_line[7][148].status_reg.re    = reg2hw.status_1940.re;


  assign rcache_line[7][149].tag_reg.tag      = reg2hw.tag_1941.q;
  assign rcache_line[7][149].tag_reg.qe       = reg2hw.tag_1941.qe;
  assign rcache_line[7][149].tag_reg.re       = reg2hw.tag_1941.re;
  assign rcache_line[7][149].status_reg.status = reg2hw.status_1941.q;//status_reg_t'(reg2hw.status_1941.q);
  assign rcache_line[7][149].status_reg.qe    = reg2hw.status_1941.qe;
  assign rcache_line[7][149].status_reg.re    = reg2hw.status_1941.re;


  assign rcache_line[7][150].tag_reg.tag      = reg2hw.tag_1942.q;
  assign rcache_line[7][150].tag_reg.qe       = reg2hw.tag_1942.qe;
  assign rcache_line[7][150].tag_reg.re       = reg2hw.tag_1942.re;
  assign rcache_line[7][150].status_reg.status = reg2hw.status_1942.q;//status_reg_t'(reg2hw.status_1942.q);
  assign rcache_line[7][150].status_reg.qe    = reg2hw.status_1942.qe;
  assign rcache_line[7][150].status_reg.re    = reg2hw.status_1942.re;


  assign rcache_line[7][151].tag_reg.tag      = reg2hw.tag_1943.q;
  assign rcache_line[7][151].tag_reg.qe       = reg2hw.tag_1943.qe;
  assign rcache_line[7][151].tag_reg.re       = reg2hw.tag_1943.re;
  assign rcache_line[7][151].status_reg.status = reg2hw.status_1943.q;//status_reg_t'(reg2hw.status_1943.q);
  assign rcache_line[7][151].status_reg.qe    = reg2hw.status_1943.qe;
  assign rcache_line[7][151].status_reg.re    = reg2hw.status_1943.re;


  assign rcache_line[7][152].tag_reg.tag      = reg2hw.tag_1944.q;
  assign rcache_line[7][152].tag_reg.qe       = reg2hw.tag_1944.qe;
  assign rcache_line[7][152].tag_reg.re       = reg2hw.tag_1944.re;
  assign rcache_line[7][152].status_reg.status = reg2hw.status_1944.q;//status_reg_t'(reg2hw.status_1944.q);
  assign rcache_line[7][152].status_reg.qe    = reg2hw.status_1944.qe;
  assign rcache_line[7][152].status_reg.re    = reg2hw.status_1944.re;


  assign rcache_line[7][153].tag_reg.tag      = reg2hw.tag_1945.q;
  assign rcache_line[7][153].tag_reg.qe       = reg2hw.tag_1945.qe;
  assign rcache_line[7][153].tag_reg.re       = reg2hw.tag_1945.re;
  assign rcache_line[7][153].status_reg.status = reg2hw.status_1945.q;//status_reg_t'(reg2hw.status_1945.q);
  assign rcache_line[7][153].status_reg.qe    = reg2hw.status_1945.qe;
  assign rcache_line[7][153].status_reg.re    = reg2hw.status_1945.re;


  assign rcache_line[7][154].tag_reg.tag      = reg2hw.tag_1946.q;
  assign rcache_line[7][154].tag_reg.qe       = reg2hw.tag_1946.qe;
  assign rcache_line[7][154].tag_reg.re       = reg2hw.tag_1946.re;
  assign rcache_line[7][154].status_reg.status = reg2hw.status_1946.q;//status_reg_t'(reg2hw.status_1946.q);
  assign rcache_line[7][154].status_reg.qe    = reg2hw.status_1946.qe;
  assign rcache_line[7][154].status_reg.re    = reg2hw.status_1946.re;


  assign rcache_line[7][155].tag_reg.tag      = reg2hw.tag_1947.q;
  assign rcache_line[7][155].tag_reg.qe       = reg2hw.tag_1947.qe;
  assign rcache_line[7][155].tag_reg.re       = reg2hw.tag_1947.re;
  assign rcache_line[7][155].status_reg.status = reg2hw.status_1947.q;//status_reg_t'(reg2hw.status_1947.q);
  assign rcache_line[7][155].status_reg.qe    = reg2hw.status_1947.qe;
  assign rcache_line[7][155].status_reg.re    = reg2hw.status_1947.re;


  assign rcache_line[7][156].tag_reg.tag      = reg2hw.tag_1948.q;
  assign rcache_line[7][156].tag_reg.qe       = reg2hw.tag_1948.qe;
  assign rcache_line[7][156].tag_reg.re       = reg2hw.tag_1948.re;
  assign rcache_line[7][156].status_reg.status = reg2hw.status_1948.q;//status_reg_t'(reg2hw.status_1948.q);
  assign rcache_line[7][156].status_reg.qe    = reg2hw.status_1948.qe;
  assign rcache_line[7][156].status_reg.re    = reg2hw.status_1948.re;


  assign rcache_line[7][157].tag_reg.tag      = reg2hw.tag_1949.q;
  assign rcache_line[7][157].tag_reg.qe       = reg2hw.tag_1949.qe;
  assign rcache_line[7][157].tag_reg.re       = reg2hw.tag_1949.re;
  assign rcache_line[7][157].status_reg.status = reg2hw.status_1949.q;//status_reg_t'(reg2hw.status_1949.q);
  assign rcache_line[7][157].status_reg.qe    = reg2hw.status_1949.qe;
  assign rcache_line[7][157].status_reg.re    = reg2hw.status_1949.re;


  assign rcache_line[7][158].tag_reg.tag      = reg2hw.tag_1950.q;
  assign rcache_line[7][158].tag_reg.qe       = reg2hw.tag_1950.qe;
  assign rcache_line[7][158].tag_reg.re       = reg2hw.tag_1950.re;
  assign rcache_line[7][158].status_reg.status = reg2hw.status_1950.q;//status_reg_t'(reg2hw.status_1950.q);
  assign rcache_line[7][158].status_reg.qe    = reg2hw.status_1950.qe;
  assign rcache_line[7][158].status_reg.re    = reg2hw.status_1950.re;


  assign rcache_line[7][159].tag_reg.tag      = reg2hw.tag_1951.q;
  assign rcache_line[7][159].tag_reg.qe       = reg2hw.tag_1951.qe;
  assign rcache_line[7][159].tag_reg.re       = reg2hw.tag_1951.re;
  assign rcache_line[7][159].status_reg.status = reg2hw.status_1951.q;//status_reg_t'(reg2hw.status_1951.q);
  assign rcache_line[7][159].status_reg.qe    = reg2hw.status_1951.qe;
  assign rcache_line[7][159].status_reg.re    = reg2hw.status_1951.re;


  assign rcache_line[7][160].tag_reg.tag      = reg2hw.tag_1952.q;
  assign rcache_line[7][160].tag_reg.qe       = reg2hw.tag_1952.qe;
  assign rcache_line[7][160].tag_reg.re       = reg2hw.tag_1952.re;
  assign rcache_line[7][160].status_reg.status = reg2hw.status_1952.q;//status_reg_t'(reg2hw.status_1952.q);
  assign rcache_line[7][160].status_reg.qe    = reg2hw.status_1952.qe;
  assign rcache_line[7][160].status_reg.re    = reg2hw.status_1952.re;


  assign rcache_line[7][161].tag_reg.tag      = reg2hw.tag_1953.q;
  assign rcache_line[7][161].tag_reg.qe       = reg2hw.tag_1953.qe;
  assign rcache_line[7][161].tag_reg.re       = reg2hw.tag_1953.re;
  assign rcache_line[7][161].status_reg.status = reg2hw.status_1953.q;//status_reg_t'(reg2hw.status_1953.q);
  assign rcache_line[7][161].status_reg.qe    = reg2hw.status_1953.qe;
  assign rcache_line[7][161].status_reg.re    = reg2hw.status_1953.re;


  assign rcache_line[7][162].tag_reg.tag      = reg2hw.tag_1954.q;
  assign rcache_line[7][162].tag_reg.qe       = reg2hw.tag_1954.qe;
  assign rcache_line[7][162].tag_reg.re       = reg2hw.tag_1954.re;
  assign rcache_line[7][162].status_reg.status = reg2hw.status_1954.q;//status_reg_t'(reg2hw.status_1954.q);
  assign rcache_line[7][162].status_reg.qe    = reg2hw.status_1954.qe;
  assign rcache_line[7][162].status_reg.re    = reg2hw.status_1954.re;


  assign rcache_line[7][163].tag_reg.tag      = reg2hw.tag_1955.q;
  assign rcache_line[7][163].tag_reg.qe       = reg2hw.tag_1955.qe;
  assign rcache_line[7][163].tag_reg.re       = reg2hw.tag_1955.re;
  assign rcache_line[7][163].status_reg.status = reg2hw.status_1955.q;//status_reg_t'(reg2hw.status_1955.q);
  assign rcache_line[7][163].status_reg.qe    = reg2hw.status_1955.qe;
  assign rcache_line[7][163].status_reg.re    = reg2hw.status_1955.re;


  assign rcache_line[7][164].tag_reg.tag      = reg2hw.tag_1956.q;
  assign rcache_line[7][164].tag_reg.qe       = reg2hw.tag_1956.qe;
  assign rcache_line[7][164].tag_reg.re       = reg2hw.tag_1956.re;
  assign rcache_line[7][164].status_reg.status = reg2hw.status_1956.q;//status_reg_t'(reg2hw.status_1956.q);
  assign rcache_line[7][164].status_reg.qe    = reg2hw.status_1956.qe;
  assign rcache_line[7][164].status_reg.re    = reg2hw.status_1956.re;


  assign rcache_line[7][165].tag_reg.tag      = reg2hw.tag_1957.q;
  assign rcache_line[7][165].tag_reg.qe       = reg2hw.tag_1957.qe;
  assign rcache_line[7][165].tag_reg.re       = reg2hw.tag_1957.re;
  assign rcache_line[7][165].status_reg.status = reg2hw.status_1957.q;//status_reg_t'(reg2hw.status_1957.q);
  assign rcache_line[7][165].status_reg.qe    = reg2hw.status_1957.qe;
  assign rcache_line[7][165].status_reg.re    = reg2hw.status_1957.re;


  assign rcache_line[7][166].tag_reg.tag      = reg2hw.tag_1958.q;
  assign rcache_line[7][166].tag_reg.qe       = reg2hw.tag_1958.qe;
  assign rcache_line[7][166].tag_reg.re       = reg2hw.tag_1958.re;
  assign rcache_line[7][166].status_reg.status = reg2hw.status_1958.q;//status_reg_t'(reg2hw.status_1958.q);
  assign rcache_line[7][166].status_reg.qe    = reg2hw.status_1958.qe;
  assign rcache_line[7][166].status_reg.re    = reg2hw.status_1958.re;


  assign rcache_line[7][167].tag_reg.tag      = reg2hw.tag_1959.q;
  assign rcache_line[7][167].tag_reg.qe       = reg2hw.tag_1959.qe;
  assign rcache_line[7][167].tag_reg.re       = reg2hw.tag_1959.re;
  assign rcache_line[7][167].status_reg.status = reg2hw.status_1959.q;//status_reg_t'(reg2hw.status_1959.q);
  assign rcache_line[7][167].status_reg.qe    = reg2hw.status_1959.qe;
  assign rcache_line[7][167].status_reg.re    = reg2hw.status_1959.re;


  assign rcache_line[7][168].tag_reg.tag      = reg2hw.tag_1960.q;
  assign rcache_line[7][168].tag_reg.qe       = reg2hw.tag_1960.qe;
  assign rcache_line[7][168].tag_reg.re       = reg2hw.tag_1960.re;
  assign rcache_line[7][168].status_reg.status = reg2hw.status_1960.q;//status_reg_t'(reg2hw.status_1960.q);
  assign rcache_line[7][168].status_reg.qe    = reg2hw.status_1960.qe;
  assign rcache_line[7][168].status_reg.re    = reg2hw.status_1960.re;


  assign rcache_line[7][169].tag_reg.tag      = reg2hw.tag_1961.q;
  assign rcache_line[7][169].tag_reg.qe       = reg2hw.tag_1961.qe;
  assign rcache_line[7][169].tag_reg.re       = reg2hw.tag_1961.re;
  assign rcache_line[7][169].status_reg.status = reg2hw.status_1961.q;//status_reg_t'(reg2hw.status_1961.q);
  assign rcache_line[7][169].status_reg.qe    = reg2hw.status_1961.qe;
  assign rcache_line[7][169].status_reg.re    = reg2hw.status_1961.re;


  assign rcache_line[7][170].tag_reg.tag      = reg2hw.tag_1962.q;
  assign rcache_line[7][170].tag_reg.qe       = reg2hw.tag_1962.qe;
  assign rcache_line[7][170].tag_reg.re       = reg2hw.tag_1962.re;
  assign rcache_line[7][170].status_reg.status = reg2hw.status_1962.q;//status_reg_t'(reg2hw.status_1962.q);
  assign rcache_line[7][170].status_reg.qe    = reg2hw.status_1962.qe;
  assign rcache_line[7][170].status_reg.re    = reg2hw.status_1962.re;


  assign rcache_line[7][171].tag_reg.tag      = reg2hw.tag_1963.q;
  assign rcache_line[7][171].tag_reg.qe       = reg2hw.tag_1963.qe;
  assign rcache_line[7][171].tag_reg.re       = reg2hw.tag_1963.re;
  assign rcache_line[7][171].status_reg.status = reg2hw.status_1963.q;//status_reg_t'(reg2hw.status_1963.q);
  assign rcache_line[7][171].status_reg.qe    = reg2hw.status_1963.qe;
  assign rcache_line[7][171].status_reg.re    = reg2hw.status_1963.re;


  assign rcache_line[7][172].tag_reg.tag      = reg2hw.tag_1964.q;
  assign rcache_line[7][172].tag_reg.qe       = reg2hw.tag_1964.qe;
  assign rcache_line[7][172].tag_reg.re       = reg2hw.tag_1964.re;
  assign rcache_line[7][172].status_reg.status = reg2hw.status_1964.q;//status_reg_t'(reg2hw.status_1964.q);
  assign rcache_line[7][172].status_reg.qe    = reg2hw.status_1964.qe;
  assign rcache_line[7][172].status_reg.re    = reg2hw.status_1964.re;


  assign rcache_line[7][173].tag_reg.tag      = reg2hw.tag_1965.q;
  assign rcache_line[7][173].tag_reg.qe       = reg2hw.tag_1965.qe;
  assign rcache_line[7][173].tag_reg.re       = reg2hw.tag_1965.re;
  assign rcache_line[7][173].status_reg.status = reg2hw.status_1965.q;//status_reg_t'(reg2hw.status_1965.q);
  assign rcache_line[7][173].status_reg.qe    = reg2hw.status_1965.qe;
  assign rcache_line[7][173].status_reg.re    = reg2hw.status_1965.re;


  assign rcache_line[7][174].tag_reg.tag      = reg2hw.tag_1966.q;
  assign rcache_line[7][174].tag_reg.qe       = reg2hw.tag_1966.qe;
  assign rcache_line[7][174].tag_reg.re       = reg2hw.tag_1966.re;
  assign rcache_line[7][174].status_reg.status = reg2hw.status_1966.q;//status_reg_t'(reg2hw.status_1966.q);
  assign rcache_line[7][174].status_reg.qe    = reg2hw.status_1966.qe;
  assign rcache_line[7][174].status_reg.re    = reg2hw.status_1966.re;


  assign rcache_line[7][175].tag_reg.tag      = reg2hw.tag_1967.q;
  assign rcache_line[7][175].tag_reg.qe       = reg2hw.tag_1967.qe;
  assign rcache_line[7][175].tag_reg.re       = reg2hw.tag_1967.re;
  assign rcache_line[7][175].status_reg.status = reg2hw.status_1967.q;//status_reg_t'(reg2hw.status_1967.q);
  assign rcache_line[7][175].status_reg.qe    = reg2hw.status_1967.qe;
  assign rcache_line[7][175].status_reg.re    = reg2hw.status_1967.re;


  assign rcache_line[7][176].tag_reg.tag      = reg2hw.tag_1968.q;
  assign rcache_line[7][176].tag_reg.qe       = reg2hw.tag_1968.qe;
  assign rcache_line[7][176].tag_reg.re       = reg2hw.tag_1968.re;
  assign rcache_line[7][176].status_reg.status = reg2hw.status_1968.q;//status_reg_t'(reg2hw.status_1968.q);
  assign rcache_line[7][176].status_reg.qe    = reg2hw.status_1968.qe;
  assign rcache_line[7][176].status_reg.re    = reg2hw.status_1968.re;


  assign rcache_line[7][177].tag_reg.tag      = reg2hw.tag_1969.q;
  assign rcache_line[7][177].tag_reg.qe       = reg2hw.tag_1969.qe;
  assign rcache_line[7][177].tag_reg.re       = reg2hw.tag_1969.re;
  assign rcache_line[7][177].status_reg.status = reg2hw.status_1969.q;//status_reg_t'(reg2hw.status_1969.q);
  assign rcache_line[7][177].status_reg.qe    = reg2hw.status_1969.qe;
  assign rcache_line[7][177].status_reg.re    = reg2hw.status_1969.re;


  assign rcache_line[7][178].tag_reg.tag      = reg2hw.tag_1970.q;
  assign rcache_line[7][178].tag_reg.qe       = reg2hw.tag_1970.qe;
  assign rcache_line[7][178].tag_reg.re       = reg2hw.tag_1970.re;
  assign rcache_line[7][178].status_reg.status = reg2hw.status_1970.q;//status_reg_t'(reg2hw.status_1970.q);
  assign rcache_line[7][178].status_reg.qe    = reg2hw.status_1970.qe;
  assign rcache_line[7][178].status_reg.re    = reg2hw.status_1970.re;


  assign rcache_line[7][179].tag_reg.tag      = reg2hw.tag_1971.q;
  assign rcache_line[7][179].tag_reg.qe       = reg2hw.tag_1971.qe;
  assign rcache_line[7][179].tag_reg.re       = reg2hw.tag_1971.re;
  assign rcache_line[7][179].status_reg.status = reg2hw.status_1971.q;//status_reg_t'(reg2hw.status_1971.q);
  assign rcache_line[7][179].status_reg.qe    = reg2hw.status_1971.qe;
  assign rcache_line[7][179].status_reg.re    = reg2hw.status_1971.re;


  assign rcache_line[7][180].tag_reg.tag      = reg2hw.tag_1972.q;
  assign rcache_line[7][180].tag_reg.qe       = reg2hw.tag_1972.qe;
  assign rcache_line[7][180].tag_reg.re       = reg2hw.tag_1972.re;
  assign rcache_line[7][180].status_reg.status = reg2hw.status_1972.q;//status_reg_t'(reg2hw.status_1972.q);
  assign rcache_line[7][180].status_reg.qe    = reg2hw.status_1972.qe;
  assign rcache_line[7][180].status_reg.re    = reg2hw.status_1972.re;


  assign rcache_line[7][181].tag_reg.tag      = reg2hw.tag_1973.q;
  assign rcache_line[7][181].tag_reg.qe       = reg2hw.tag_1973.qe;
  assign rcache_line[7][181].tag_reg.re       = reg2hw.tag_1973.re;
  assign rcache_line[7][181].status_reg.status = reg2hw.status_1973.q;//status_reg_t'(reg2hw.status_1973.q);
  assign rcache_line[7][181].status_reg.qe    = reg2hw.status_1973.qe;
  assign rcache_line[7][181].status_reg.re    = reg2hw.status_1973.re;


  assign rcache_line[7][182].tag_reg.tag      = reg2hw.tag_1974.q;
  assign rcache_line[7][182].tag_reg.qe       = reg2hw.tag_1974.qe;
  assign rcache_line[7][182].tag_reg.re       = reg2hw.tag_1974.re;
  assign rcache_line[7][182].status_reg.status = reg2hw.status_1974.q;//status_reg_t'(reg2hw.status_1974.q);
  assign rcache_line[7][182].status_reg.qe    = reg2hw.status_1974.qe;
  assign rcache_line[7][182].status_reg.re    = reg2hw.status_1974.re;


  assign rcache_line[7][183].tag_reg.tag      = reg2hw.tag_1975.q;
  assign rcache_line[7][183].tag_reg.qe       = reg2hw.tag_1975.qe;
  assign rcache_line[7][183].tag_reg.re       = reg2hw.tag_1975.re;
  assign rcache_line[7][183].status_reg.status = reg2hw.status_1975.q;//status_reg_t'(reg2hw.status_1975.q);
  assign rcache_line[7][183].status_reg.qe    = reg2hw.status_1975.qe;
  assign rcache_line[7][183].status_reg.re    = reg2hw.status_1975.re;


  assign rcache_line[7][184].tag_reg.tag      = reg2hw.tag_1976.q;
  assign rcache_line[7][184].tag_reg.qe       = reg2hw.tag_1976.qe;
  assign rcache_line[7][184].tag_reg.re       = reg2hw.tag_1976.re;
  assign rcache_line[7][184].status_reg.status = reg2hw.status_1976.q;//status_reg_t'(reg2hw.status_1976.q);
  assign rcache_line[7][184].status_reg.qe    = reg2hw.status_1976.qe;
  assign rcache_line[7][184].status_reg.re    = reg2hw.status_1976.re;


  assign rcache_line[7][185].tag_reg.tag      = reg2hw.tag_1977.q;
  assign rcache_line[7][185].tag_reg.qe       = reg2hw.tag_1977.qe;
  assign rcache_line[7][185].tag_reg.re       = reg2hw.tag_1977.re;
  assign rcache_line[7][185].status_reg.status = reg2hw.status_1977.q;//status_reg_t'(reg2hw.status_1977.q);
  assign rcache_line[7][185].status_reg.qe    = reg2hw.status_1977.qe;
  assign rcache_line[7][185].status_reg.re    = reg2hw.status_1977.re;


  assign rcache_line[7][186].tag_reg.tag      = reg2hw.tag_1978.q;
  assign rcache_line[7][186].tag_reg.qe       = reg2hw.tag_1978.qe;
  assign rcache_line[7][186].tag_reg.re       = reg2hw.tag_1978.re;
  assign rcache_line[7][186].status_reg.status = reg2hw.status_1978.q;//status_reg_t'(reg2hw.status_1978.q);
  assign rcache_line[7][186].status_reg.qe    = reg2hw.status_1978.qe;
  assign rcache_line[7][186].status_reg.re    = reg2hw.status_1978.re;


  assign rcache_line[7][187].tag_reg.tag      = reg2hw.tag_1979.q;
  assign rcache_line[7][187].tag_reg.qe       = reg2hw.tag_1979.qe;
  assign rcache_line[7][187].tag_reg.re       = reg2hw.tag_1979.re;
  assign rcache_line[7][187].status_reg.status = reg2hw.status_1979.q;//status_reg_t'(reg2hw.status_1979.q);
  assign rcache_line[7][187].status_reg.qe    = reg2hw.status_1979.qe;
  assign rcache_line[7][187].status_reg.re    = reg2hw.status_1979.re;


  assign rcache_line[7][188].tag_reg.tag      = reg2hw.tag_1980.q;
  assign rcache_line[7][188].tag_reg.qe       = reg2hw.tag_1980.qe;
  assign rcache_line[7][188].tag_reg.re       = reg2hw.tag_1980.re;
  assign rcache_line[7][188].status_reg.status = reg2hw.status_1980.q;//status_reg_t'(reg2hw.status_1980.q);
  assign rcache_line[7][188].status_reg.qe    = reg2hw.status_1980.qe;
  assign rcache_line[7][188].status_reg.re    = reg2hw.status_1980.re;


  assign rcache_line[7][189].tag_reg.tag      = reg2hw.tag_1981.q;
  assign rcache_line[7][189].tag_reg.qe       = reg2hw.tag_1981.qe;
  assign rcache_line[7][189].tag_reg.re       = reg2hw.tag_1981.re;
  assign rcache_line[7][189].status_reg.status = reg2hw.status_1981.q;//status_reg_t'(reg2hw.status_1981.q);
  assign rcache_line[7][189].status_reg.qe    = reg2hw.status_1981.qe;
  assign rcache_line[7][189].status_reg.re    = reg2hw.status_1981.re;


  assign rcache_line[7][190].tag_reg.tag      = reg2hw.tag_1982.q;
  assign rcache_line[7][190].tag_reg.qe       = reg2hw.tag_1982.qe;
  assign rcache_line[7][190].tag_reg.re       = reg2hw.tag_1982.re;
  assign rcache_line[7][190].status_reg.status = reg2hw.status_1982.q;//status_reg_t'(reg2hw.status_1982.q);
  assign rcache_line[7][190].status_reg.qe    = reg2hw.status_1982.qe;
  assign rcache_line[7][190].status_reg.re    = reg2hw.status_1982.re;


  assign rcache_line[7][191].tag_reg.tag      = reg2hw.tag_1983.q;
  assign rcache_line[7][191].tag_reg.qe       = reg2hw.tag_1983.qe;
  assign rcache_line[7][191].tag_reg.re       = reg2hw.tag_1983.re;
  assign rcache_line[7][191].status_reg.status = reg2hw.status_1983.q;//status_reg_t'(reg2hw.status_1983.q);
  assign rcache_line[7][191].status_reg.qe    = reg2hw.status_1983.qe;
  assign rcache_line[7][191].status_reg.re    = reg2hw.status_1983.re;


  assign rcache_line[7][192].tag_reg.tag      = reg2hw.tag_1984.q;
  assign rcache_line[7][192].tag_reg.qe       = reg2hw.tag_1984.qe;
  assign rcache_line[7][192].tag_reg.re       = reg2hw.tag_1984.re;
  assign rcache_line[7][192].status_reg.status = reg2hw.status_1984.q;//status_reg_t'(reg2hw.status_1984.q);
  assign rcache_line[7][192].status_reg.qe    = reg2hw.status_1984.qe;
  assign rcache_line[7][192].status_reg.re    = reg2hw.status_1984.re;


  assign rcache_line[7][193].tag_reg.tag      = reg2hw.tag_1985.q;
  assign rcache_line[7][193].tag_reg.qe       = reg2hw.tag_1985.qe;
  assign rcache_line[7][193].tag_reg.re       = reg2hw.tag_1985.re;
  assign rcache_line[7][193].status_reg.status = reg2hw.status_1985.q;//status_reg_t'(reg2hw.status_1985.q);
  assign rcache_line[7][193].status_reg.qe    = reg2hw.status_1985.qe;
  assign rcache_line[7][193].status_reg.re    = reg2hw.status_1985.re;


  assign rcache_line[7][194].tag_reg.tag      = reg2hw.tag_1986.q;
  assign rcache_line[7][194].tag_reg.qe       = reg2hw.tag_1986.qe;
  assign rcache_line[7][194].tag_reg.re       = reg2hw.tag_1986.re;
  assign rcache_line[7][194].status_reg.status = reg2hw.status_1986.q;//status_reg_t'(reg2hw.status_1986.q);
  assign rcache_line[7][194].status_reg.qe    = reg2hw.status_1986.qe;
  assign rcache_line[7][194].status_reg.re    = reg2hw.status_1986.re;


  assign rcache_line[7][195].tag_reg.tag      = reg2hw.tag_1987.q;
  assign rcache_line[7][195].tag_reg.qe       = reg2hw.tag_1987.qe;
  assign rcache_line[7][195].tag_reg.re       = reg2hw.tag_1987.re;
  assign rcache_line[7][195].status_reg.status = reg2hw.status_1987.q;//status_reg_t'(reg2hw.status_1987.q);
  assign rcache_line[7][195].status_reg.qe    = reg2hw.status_1987.qe;
  assign rcache_line[7][195].status_reg.re    = reg2hw.status_1987.re;


  assign rcache_line[7][196].tag_reg.tag      = reg2hw.tag_1988.q;
  assign rcache_line[7][196].tag_reg.qe       = reg2hw.tag_1988.qe;
  assign rcache_line[7][196].tag_reg.re       = reg2hw.tag_1988.re;
  assign rcache_line[7][196].status_reg.status = reg2hw.status_1988.q;//status_reg_t'(reg2hw.status_1988.q);
  assign rcache_line[7][196].status_reg.qe    = reg2hw.status_1988.qe;
  assign rcache_line[7][196].status_reg.re    = reg2hw.status_1988.re;


  assign rcache_line[7][197].tag_reg.tag      = reg2hw.tag_1989.q;
  assign rcache_line[7][197].tag_reg.qe       = reg2hw.tag_1989.qe;
  assign rcache_line[7][197].tag_reg.re       = reg2hw.tag_1989.re;
  assign rcache_line[7][197].status_reg.status = reg2hw.status_1989.q;//status_reg_t'(reg2hw.status_1989.q);
  assign rcache_line[7][197].status_reg.qe    = reg2hw.status_1989.qe;
  assign rcache_line[7][197].status_reg.re    = reg2hw.status_1989.re;


  assign rcache_line[7][198].tag_reg.tag      = reg2hw.tag_1990.q;
  assign rcache_line[7][198].tag_reg.qe       = reg2hw.tag_1990.qe;
  assign rcache_line[7][198].tag_reg.re       = reg2hw.tag_1990.re;
  assign rcache_line[7][198].status_reg.status = reg2hw.status_1990.q;//status_reg_t'(reg2hw.status_1990.q);
  assign rcache_line[7][198].status_reg.qe    = reg2hw.status_1990.qe;
  assign rcache_line[7][198].status_reg.re    = reg2hw.status_1990.re;


  assign rcache_line[7][199].tag_reg.tag      = reg2hw.tag_1991.q;
  assign rcache_line[7][199].tag_reg.qe       = reg2hw.tag_1991.qe;
  assign rcache_line[7][199].tag_reg.re       = reg2hw.tag_1991.re;
  assign rcache_line[7][199].status_reg.status = reg2hw.status_1991.q;//status_reg_t'(reg2hw.status_1991.q);
  assign rcache_line[7][199].status_reg.qe    = reg2hw.status_1991.qe;
  assign rcache_line[7][199].status_reg.re    = reg2hw.status_1991.re;


  assign rcache_line[7][200].tag_reg.tag      = reg2hw.tag_1992.q;
  assign rcache_line[7][200].tag_reg.qe       = reg2hw.tag_1992.qe;
  assign rcache_line[7][200].tag_reg.re       = reg2hw.tag_1992.re;
  assign rcache_line[7][200].status_reg.status = reg2hw.status_1992.q;//status_reg_t'(reg2hw.status_1992.q);
  assign rcache_line[7][200].status_reg.qe    = reg2hw.status_1992.qe;
  assign rcache_line[7][200].status_reg.re    = reg2hw.status_1992.re;


  assign rcache_line[7][201].tag_reg.tag      = reg2hw.tag_1993.q;
  assign rcache_line[7][201].tag_reg.qe       = reg2hw.tag_1993.qe;
  assign rcache_line[7][201].tag_reg.re       = reg2hw.tag_1993.re;
  assign rcache_line[7][201].status_reg.status = reg2hw.status_1993.q;//status_reg_t'(reg2hw.status_1993.q);
  assign rcache_line[7][201].status_reg.qe    = reg2hw.status_1993.qe;
  assign rcache_line[7][201].status_reg.re    = reg2hw.status_1993.re;


  assign rcache_line[7][202].tag_reg.tag      = reg2hw.tag_1994.q;
  assign rcache_line[7][202].tag_reg.qe       = reg2hw.tag_1994.qe;
  assign rcache_line[7][202].tag_reg.re       = reg2hw.tag_1994.re;
  assign rcache_line[7][202].status_reg.status = reg2hw.status_1994.q;//status_reg_t'(reg2hw.status_1994.q);
  assign rcache_line[7][202].status_reg.qe    = reg2hw.status_1994.qe;
  assign rcache_line[7][202].status_reg.re    = reg2hw.status_1994.re;


  assign rcache_line[7][203].tag_reg.tag      = reg2hw.tag_1995.q;
  assign rcache_line[7][203].tag_reg.qe       = reg2hw.tag_1995.qe;
  assign rcache_line[7][203].tag_reg.re       = reg2hw.tag_1995.re;
  assign rcache_line[7][203].status_reg.status = reg2hw.status_1995.q;//status_reg_t'(reg2hw.status_1995.q);
  assign rcache_line[7][203].status_reg.qe    = reg2hw.status_1995.qe;
  assign rcache_line[7][203].status_reg.re    = reg2hw.status_1995.re;


  assign rcache_line[7][204].tag_reg.tag      = reg2hw.tag_1996.q;
  assign rcache_line[7][204].tag_reg.qe       = reg2hw.tag_1996.qe;
  assign rcache_line[7][204].tag_reg.re       = reg2hw.tag_1996.re;
  assign rcache_line[7][204].status_reg.status = reg2hw.status_1996.q;//status_reg_t'(reg2hw.status_1996.q);
  assign rcache_line[7][204].status_reg.qe    = reg2hw.status_1996.qe;
  assign rcache_line[7][204].status_reg.re    = reg2hw.status_1996.re;


  assign rcache_line[7][205].tag_reg.tag      = reg2hw.tag_1997.q;
  assign rcache_line[7][205].tag_reg.qe       = reg2hw.tag_1997.qe;
  assign rcache_line[7][205].tag_reg.re       = reg2hw.tag_1997.re;
  assign rcache_line[7][205].status_reg.status = reg2hw.status_1997.q;//status_reg_t'(reg2hw.status_1997.q);
  assign rcache_line[7][205].status_reg.qe    = reg2hw.status_1997.qe;
  assign rcache_line[7][205].status_reg.re    = reg2hw.status_1997.re;


  assign rcache_line[7][206].tag_reg.tag      = reg2hw.tag_1998.q;
  assign rcache_line[7][206].tag_reg.qe       = reg2hw.tag_1998.qe;
  assign rcache_line[7][206].tag_reg.re       = reg2hw.tag_1998.re;
  assign rcache_line[7][206].status_reg.status = reg2hw.status_1998.q;//status_reg_t'(reg2hw.status_1998.q);
  assign rcache_line[7][206].status_reg.qe    = reg2hw.status_1998.qe;
  assign rcache_line[7][206].status_reg.re    = reg2hw.status_1998.re;


  assign rcache_line[7][207].tag_reg.tag      = reg2hw.tag_1999.q;
  assign rcache_line[7][207].tag_reg.qe       = reg2hw.tag_1999.qe;
  assign rcache_line[7][207].tag_reg.re       = reg2hw.tag_1999.re;
  assign rcache_line[7][207].status_reg.status = reg2hw.status_1999.q;//status_reg_t'(reg2hw.status_1999.q);
  assign rcache_line[7][207].status_reg.qe    = reg2hw.status_1999.qe;
  assign rcache_line[7][207].status_reg.re    = reg2hw.status_1999.re;


  assign rcache_line[7][208].tag_reg.tag      = reg2hw.tag_2000.q;
  assign rcache_line[7][208].tag_reg.qe       = reg2hw.tag_2000.qe;
  assign rcache_line[7][208].tag_reg.re       = reg2hw.tag_2000.re;
  assign rcache_line[7][208].status_reg.status = reg2hw.status_2000.q;//status_reg_t'(reg2hw.status_2000.q);
  assign rcache_line[7][208].status_reg.qe    = reg2hw.status_2000.qe;
  assign rcache_line[7][208].status_reg.re    = reg2hw.status_2000.re;


  assign rcache_line[7][209].tag_reg.tag      = reg2hw.tag_2001.q;
  assign rcache_line[7][209].tag_reg.qe       = reg2hw.tag_2001.qe;
  assign rcache_line[7][209].tag_reg.re       = reg2hw.tag_2001.re;
  assign rcache_line[7][209].status_reg.status = reg2hw.status_2001.q;//status_reg_t'(reg2hw.status_2001.q);
  assign rcache_line[7][209].status_reg.qe    = reg2hw.status_2001.qe;
  assign rcache_line[7][209].status_reg.re    = reg2hw.status_2001.re;


  assign rcache_line[7][210].tag_reg.tag      = reg2hw.tag_2002.q;
  assign rcache_line[7][210].tag_reg.qe       = reg2hw.tag_2002.qe;
  assign rcache_line[7][210].tag_reg.re       = reg2hw.tag_2002.re;
  assign rcache_line[7][210].status_reg.status = reg2hw.status_2002.q;//status_reg_t'(reg2hw.status_2002.q);
  assign rcache_line[7][210].status_reg.qe    = reg2hw.status_2002.qe;
  assign rcache_line[7][210].status_reg.re    = reg2hw.status_2002.re;


  assign rcache_line[7][211].tag_reg.tag      = reg2hw.tag_2003.q;
  assign rcache_line[7][211].tag_reg.qe       = reg2hw.tag_2003.qe;
  assign rcache_line[7][211].tag_reg.re       = reg2hw.tag_2003.re;
  assign rcache_line[7][211].status_reg.status = reg2hw.status_2003.q;//status_reg_t'(reg2hw.status_2003.q);
  assign rcache_line[7][211].status_reg.qe    = reg2hw.status_2003.qe;
  assign rcache_line[7][211].status_reg.re    = reg2hw.status_2003.re;


  assign rcache_line[7][212].tag_reg.tag      = reg2hw.tag_2004.q;
  assign rcache_line[7][212].tag_reg.qe       = reg2hw.tag_2004.qe;
  assign rcache_line[7][212].tag_reg.re       = reg2hw.tag_2004.re;
  assign rcache_line[7][212].status_reg.status = reg2hw.status_2004.q;//status_reg_t'(reg2hw.status_2004.q);
  assign rcache_line[7][212].status_reg.qe    = reg2hw.status_2004.qe;
  assign rcache_line[7][212].status_reg.re    = reg2hw.status_2004.re;


  assign rcache_line[7][213].tag_reg.tag      = reg2hw.tag_2005.q;
  assign rcache_line[7][213].tag_reg.qe       = reg2hw.tag_2005.qe;
  assign rcache_line[7][213].tag_reg.re       = reg2hw.tag_2005.re;
  assign rcache_line[7][213].status_reg.status = reg2hw.status_2005.q;//status_reg_t'(reg2hw.status_2005.q);
  assign rcache_line[7][213].status_reg.qe    = reg2hw.status_2005.qe;
  assign rcache_line[7][213].status_reg.re    = reg2hw.status_2005.re;


  assign rcache_line[7][214].tag_reg.tag      = reg2hw.tag_2006.q;
  assign rcache_line[7][214].tag_reg.qe       = reg2hw.tag_2006.qe;
  assign rcache_line[7][214].tag_reg.re       = reg2hw.tag_2006.re;
  assign rcache_line[7][214].status_reg.status = reg2hw.status_2006.q;//status_reg_t'(reg2hw.status_2006.q);
  assign rcache_line[7][214].status_reg.qe    = reg2hw.status_2006.qe;
  assign rcache_line[7][214].status_reg.re    = reg2hw.status_2006.re;


  assign rcache_line[7][215].tag_reg.tag      = reg2hw.tag_2007.q;
  assign rcache_line[7][215].tag_reg.qe       = reg2hw.tag_2007.qe;
  assign rcache_line[7][215].tag_reg.re       = reg2hw.tag_2007.re;
  assign rcache_line[7][215].status_reg.status = reg2hw.status_2007.q;//status_reg_t'(reg2hw.status_2007.q);
  assign rcache_line[7][215].status_reg.qe    = reg2hw.status_2007.qe;
  assign rcache_line[7][215].status_reg.re    = reg2hw.status_2007.re;


  assign rcache_line[7][216].tag_reg.tag      = reg2hw.tag_2008.q;
  assign rcache_line[7][216].tag_reg.qe       = reg2hw.tag_2008.qe;
  assign rcache_line[7][216].tag_reg.re       = reg2hw.tag_2008.re;
  assign rcache_line[7][216].status_reg.status = reg2hw.status_2008.q;//status_reg_t'(reg2hw.status_2008.q);
  assign rcache_line[7][216].status_reg.qe    = reg2hw.status_2008.qe;
  assign rcache_line[7][216].status_reg.re    = reg2hw.status_2008.re;


  assign rcache_line[7][217].tag_reg.tag      = reg2hw.tag_2009.q;
  assign rcache_line[7][217].tag_reg.qe       = reg2hw.tag_2009.qe;
  assign rcache_line[7][217].tag_reg.re       = reg2hw.tag_2009.re;
  assign rcache_line[7][217].status_reg.status = reg2hw.status_2009.q;//status_reg_t'(reg2hw.status_2009.q);
  assign rcache_line[7][217].status_reg.qe    = reg2hw.status_2009.qe;
  assign rcache_line[7][217].status_reg.re    = reg2hw.status_2009.re;


  assign rcache_line[7][218].tag_reg.tag      = reg2hw.tag_2010.q;
  assign rcache_line[7][218].tag_reg.qe       = reg2hw.tag_2010.qe;
  assign rcache_line[7][218].tag_reg.re       = reg2hw.tag_2010.re;
  assign rcache_line[7][218].status_reg.status = reg2hw.status_2010.q;//status_reg_t'(reg2hw.status_2010.q);
  assign rcache_line[7][218].status_reg.qe    = reg2hw.status_2010.qe;
  assign rcache_line[7][218].status_reg.re    = reg2hw.status_2010.re;


  assign rcache_line[7][219].tag_reg.tag      = reg2hw.tag_2011.q;
  assign rcache_line[7][219].tag_reg.qe       = reg2hw.tag_2011.qe;
  assign rcache_line[7][219].tag_reg.re       = reg2hw.tag_2011.re;
  assign rcache_line[7][219].status_reg.status = reg2hw.status_2011.q;//status_reg_t'(reg2hw.status_2011.q);
  assign rcache_line[7][219].status_reg.qe    = reg2hw.status_2011.qe;
  assign rcache_line[7][219].status_reg.re    = reg2hw.status_2011.re;


  assign rcache_line[7][220].tag_reg.tag      = reg2hw.tag_2012.q;
  assign rcache_line[7][220].tag_reg.qe       = reg2hw.tag_2012.qe;
  assign rcache_line[7][220].tag_reg.re       = reg2hw.tag_2012.re;
  assign rcache_line[7][220].status_reg.status = reg2hw.status_2012.q;//status_reg_t'(reg2hw.status_2012.q);
  assign rcache_line[7][220].status_reg.qe    = reg2hw.status_2012.qe;
  assign rcache_line[7][220].status_reg.re    = reg2hw.status_2012.re;


  assign rcache_line[7][221].tag_reg.tag      = reg2hw.tag_2013.q;
  assign rcache_line[7][221].tag_reg.qe       = reg2hw.tag_2013.qe;
  assign rcache_line[7][221].tag_reg.re       = reg2hw.tag_2013.re;
  assign rcache_line[7][221].status_reg.status = reg2hw.status_2013.q;//status_reg_t'(reg2hw.status_2013.q);
  assign rcache_line[7][221].status_reg.qe    = reg2hw.status_2013.qe;
  assign rcache_line[7][221].status_reg.re    = reg2hw.status_2013.re;


  assign rcache_line[7][222].tag_reg.tag      = reg2hw.tag_2014.q;
  assign rcache_line[7][222].tag_reg.qe       = reg2hw.tag_2014.qe;
  assign rcache_line[7][222].tag_reg.re       = reg2hw.tag_2014.re;
  assign rcache_line[7][222].status_reg.status = reg2hw.status_2014.q;//status_reg_t'(reg2hw.status_2014.q);
  assign rcache_line[7][222].status_reg.qe    = reg2hw.status_2014.qe;
  assign rcache_line[7][222].status_reg.re    = reg2hw.status_2014.re;


  assign rcache_line[7][223].tag_reg.tag      = reg2hw.tag_2015.q;
  assign rcache_line[7][223].tag_reg.qe       = reg2hw.tag_2015.qe;
  assign rcache_line[7][223].tag_reg.re       = reg2hw.tag_2015.re;
  assign rcache_line[7][223].status_reg.status = reg2hw.status_2015.q;//status_reg_t'(reg2hw.status_2015.q);
  assign rcache_line[7][223].status_reg.qe    = reg2hw.status_2015.qe;
  assign rcache_line[7][223].status_reg.re    = reg2hw.status_2015.re;


  assign rcache_line[7][224].tag_reg.tag      = reg2hw.tag_2016.q;
  assign rcache_line[7][224].tag_reg.qe       = reg2hw.tag_2016.qe;
  assign rcache_line[7][224].tag_reg.re       = reg2hw.tag_2016.re;
  assign rcache_line[7][224].status_reg.status = reg2hw.status_2016.q;//status_reg_t'(reg2hw.status_2016.q);
  assign rcache_line[7][224].status_reg.qe    = reg2hw.status_2016.qe;
  assign rcache_line[7][224].status_reg.re    = reg2hw.status_2016.re;


  assign rcache_line[7][225].tag_reg.tag      = reg2hw.tag_2017.q;
  assign rcache_line[7][225].tag_reg.qe       = reg2hw.tag_2017.qe;
  assign rcache_line[7][225].tag_reg.re       = reg2hw.tag_2017.re;
  assign rcache_line[7][225].status_reg.status = reg2hw.status_2017.q;//status_reg_t'(reg2hw.status_2017.q);
  assign rcache_line[7][225].status_reg.qe    = reg2hw.status_2017.qe;
  assign rcache_line[7][225].status_reg.re    = reg2hw.status_2017.re;


  assign rcache_line[7][226].tag_reg.tag      = reg2hw.tag_2018.q;
  assign rcache_line[7][226].tag_reg.qe       = reg2hw.tag_2018.qe;
  assign rcache_line[7][226].tag_reg.re       = reg2hw.tag_2018.re;
  assign rcache_line[7][226].status_reg.status = reg2hw.status_2018.q;//status_reg_t'(reg2hw.status_2018.q);
  assign rcache_line[7][226].status_reg.qe    = reg2hw.status_2018.qe;
  assign rcache_line[7][226].status_reg.re    = reg2hw.status_2018.re;


  assign rcache_line[7][227].tag_reg.tag      = reg2hw.tag_2019.q;
  assign rcache_line[7][227].tag_reg.qe       = reg2hw.tag_2019.qe;
  assign rcache_line[7][227].tag_reg.re       = reg2hw.tag_2019.re;
  assign rcache_line[7][227].status_reg.status = reg2hw.status_2019.q;//status_reg_t'(reg2hw.status_2019.q);
  assign rcache_line[7][227].status_reg.qe    = reg2hw.status_2019.qe;
  assign rcache_line[7][227].status_reg.re    = reg2hw.status_2019.re;


  assign rcache_line[7][228].tag_reg.tag      = reg2hw.tag_2020.q;
  assign rcache_line[7][228].tag_reg.qe       = reg2hw.tag_2020.qe;
  assign rcache_line[7][228].tag_reg.re       = reg2hw.tag_2020.re;
  assign rcache_line[7][228].status_reg.status = reg2hw.status_2020.q;//status_reg_t'(reg2hw.status_2020.q);
  assign rcache_line[7][228].status_reg.qe    = reg2hw.status_2020.qe;
  assign rcache_line[7][228].status_reg.re    = reg2hw.status_2020.re;


  assign rcache_line[7][229].tag_reg.tag      = reg2hw.tag_2021.q;
  assign rcache_line[7][229].tag_reg.qe       = reg2hw.tag_2021.qe;
  assign rcache_line[7][229].tag_reg.re       = reg2hw.tag_2021.re;
  assign rcache_line[7][229].status_reg.status = reg2hw.status_2021.q;//status_reg_t'(reg2hw.status_2021.q);
  assign rcache_line[7][229].status_reg.qe    = reg2hw.status_2021.qe;
  assign rcache_line[7][229].status_reg.re    = reg2hw.status_2021.re;


  assign rcache_line[7][230].tag_reg.tag      = reg2hw.tag_2022.q;
  assign rcache_line[7][230].tag_reg.qe       = reg2hw.tag_2022.qe;
  assign rcache_line[7][230].tag_reg.re       = reg2hw.tag_2022.re;
  assign rcache_line[7][230].status_reg.status = reg2hw.status_2022.q;//status_reg_t'(reg2hw.status_2022.q);
  assign rcache_line[7][230].status_reg.qe    = reg2hw.status_2022.qe;
  assign rcache_line[7][230].status_reg.re    = reg2hw.status_2022.re;


  assign rcache_line[7][231].tag_reg.tag      = reg2hw.tag_2023.q;
  assign rcache_line[7][231].tag_reg.qe       = reg2hw.tag_2023.qe;
  assign rcache_line[7][231].tag_reg.re       = reg2hw.tag_2023.re;
  assign rcache_line[7][231].status_reg.status = reg2hw.status_2023.q;//status_reg_t'(reg2hw.status_2023.q);
  assign rcache_line[7][231].status_reg.qe    = reg2hw.status_2023.qe;
  assign rcache_line[7][231].status_reg.re    = reg2hw.status_2023.re;


  assign rcache_line[7][232].tag_reg.tag      = reg2hw.tag_2024.q;
  assign rcache_line[7][232].tag_reg.qe       = reg2hw.tag_2024.qe;
  assign rcache_line[7][232].tag_reg.re       = reg2hw.tag_2024.re;
  assign rcache_line[7][232].status_reg.status = reg2hw.status_2024.q;//status_reg_t'(reg2hw.status_2024.q);
  assign rcache_line[7][232].status_reg.qe    = reg2hw.status_2024.qe;
  assign rcache_line[7][232].status_reg.re    = reg2hw.status_2024.re;


  assign rcache_line[7][233].tag_reg.tag      = reg2hw.tag_2025.q;
  assign rcache_line[7][233].tag_reg.qe       = reg2hw.tag_2025.qe;
  assign rcache_line[7][233].tag_reg.re       = reg2hw.tag_2025.re;
  assign rcache_line[7][233].status_reg.status = reg2hw.status_2025.q;//status_reg_t'(reg2hw.status_2025.q);
  assign rcache_line[7][233].status_reg.qe    = reg2hw.status_2025.qe;
  assign rcache_line[7][233].status_reg.re    = reg2hw.status_2025.re;


  assign rcache_line[7][234].tag_reg.tag      = reg2hw.tag_2026.q;
  assign rcache_line[7][234].tag_reg.qe       = reg2hw.tag_2026.qe;
  assign rcache_line[7][234].tag_reg.re       = reg2hw.tag_2026.re;
  assign rcache_line[7][234].status_reg.status = reg2hw.status_2026.q;//status_reg_t'(reg2hw.status_2026.q);
  assign rcache_line[7][234].status_reg.qe    = reg2hw.status_2026.qe;
  assign rcache_line[7][234].status_reg.re    = reg2hw.status_2026.re;


  assign rcache_line[7][235].tag_reg.tag      = reg2hw.tag_2027.q;
  assign rcache_line[7][235].tag_reg.qe       = reg2hw.tag_2027.qe;
  assign rcache_line[7][235].tag_reg.re       = reg2hw.tag_2027.re;
  assign rcache_line[7][235].status_reg.status = reg2hw.status_2027.q;//status_reg_t'(reg2hw.status_2027.q);
  assign rcache_line[7][235].status_reg.qe    = reg2hw.status_2027.qe;
  assign rcache_line[7][235].status_reg.re    = reg2hw.status_2027.re;


  assign rcache_line[7][236].tag_reg.tag      = reg2hw.tag_2028.q;
  assign rcache_line[7][236].tag_reg.qe       = reg2hw.tag_2028.qe;
  assign rcache_line[7][236].tag_reg.re       = reg2hw.tag_2028.re;
  assign rcache_line[7][236].status_reg.status = reg2hw.status_2028.q;//status_reg_t'(reg2hw.status_2028.q);
  assign rcache_line[7][236].status_reg.qe    = reg2hw.status_2028.qe;
  assign rcache_line[7][236].status_reg.re    = reg2hw.status_2028.re;


  assign rcache_line[7][237].tag_reg.tag      = reg2hw.tag_2029.q;
  assign rcache_line[7][237].tag_reg.qe       = reg2hw.tag_2029.qe;
  assign rcache_line[7][237].tag_reg.re       = reg2hw.tag_2029.re;
  assign rcache_line[7][237].status_reg.status = reg2hw.status_2029.q;//status_reg_t'(reg2hw.status_2029.q);
  assign rcache_line[7][237].status_reg.qe    = reg2hw.status_2029.qe;
  assign rcache_line[7][237].status_reg.re    = reg2hw.status_2029.re;


  assign rcache_line[7][238].tag_reg.tag      = reg2hw.tag_2030.q;
  assign rcache_line[7][238].tag_reg.qe       = reg2hw.tag_2030.qe;
  assign rcache_line[7][238].tag_reg.re       = reg2hw.tag_2030.re;
  assign rcache_line[7][238].status_reg.status = reg2hw.status_2030.q;//status_reg_t'(reg2hw.status_2030.q);
  assign rcache_line[7][238].status_reg.qe    = reg2hw.status_2030.qe;
  assign rcache_line[7][238].status_reg.re    = reg2hw.status_2030.re;


  assign rcache_line[7][239].tag_reg.tag      = reg2hw.tag_2031.q;
  assign rcache_line[7][239].tag_reg.qe       = reg2hw.tag_2031.qe;
  assign rcache_line[7][239].tag_reg.re       = reg2hw.tag_2031.re;
  assign rcache_line[7][239].status_reg.status = reg2hw.status_2031.q;//status_reg_t'(reg2hw.status_2031.q);
  assign rcache_line[7][239].status_reg.qe    = reg2hw.status_2031.qe;
  assign rcache_line[7][239].status_reg.re    = reg2hw.status_2031.re;


  assign rcache_line[7][240].tag_reg.tag      = reg2hw.tag_2032.q;
  assign rcache_line[7][240].tag_reg.qe       = reg2hw.tag_2032.qe;
  assign rcache_line[7][240].tag_reg.re       = reg2hw.tag_2032.re;
  assign rcache_line[7][240].status_reg.status = reg2hw.status_2032.q;//status_reg_t'(reg2hw.status_2032.q);
  assign rcache_line[7][240].status_reg.qe    = reg2hw.status_2032.qe;
  assign rcache_line[7][240].status_reg.re    = reg2hw.status_2032.re;


  assign rcache_line[7][241].tag_reg.tag      = reg2hw.tag_2033.q;
  assign rcache_line[7][241].tag_reg.qe       = reg2hw.tag_2033.qe;
  assign rcache_line[7][241].tag_reg.re       = reg2hw.tag_2033.re;
  assign rcache_line[7][241].status_reg.status = reg2hw.status_2033.q;//status_reg_t'(reg2hw.status_2033.q);
  assign rcache_line[7][241].status_reg.qe    = reg2hw.status_2033.qe;
  assign rcache_line[7][241].status_reg.re    = reg2hw.status_2033.re;


  assign rcache_line[7][242].tag_reg.tag      = reg2hw.tag_2034.q;
  assign rcache_line[7][242].tag_reg.qe       = reg2hw.tag_2034.qe;
  assign rcache_line[7][242].tag_reg.re       = reg2hw.tag_2034.re;
  assign rcache_line[7][242].status_reg.status = reg2hw.status_2034.q;//status_reg_t'(reg2hw.status_2034.q);
  assign rcache_line[7][242].status_reg.qe    = reg2hw.status_2034.qe;
  assign rcache_line[7][242].status_reg.re    = reg2hw.status_2034.re;


  assign rcache_line[7][243].tag_reg.tag      = reg2hw.tag_2035.q;
  assign rcache_line[7][243].tag_reg.qe       = reg2hw.tag_2035.qe;
  assign rcache_line[7][243].tag_reg.re       = reg2hw.tag_2035.re;
  assign rcache_line[7][243].status_reg.status = reg2hw.status_2035.q;//status_reg_t'(reg2hw.status_2035.q);
  assign rcache_line[7][243].status_reg.qe    = reg2hw.status_2035.qe;
  assign rcache_line[7][243].status_reg.re    = reg2hw.status_2035.re;


  assign rcache_line[7][244].tag_reg.tag      = reg2hw.tag_2036.q;
  assign rcache_line[7][244].tag_reg.qe       = reg2hw.tag_2036.qe;
  assign rcache_line[7][244].tag_reg.re       = reg2hw.tag_2036.re;
  assign rcache_line[7][244].status_reg.status = reg2hw.status_2036.q;//status_reg_t'(reg2hw.status_2036.q);
  assign rcache_line[7][244].status_reg.qe    = reg2hw.status_2036.qe;
  assign rcache_line[7][244].status_reg.re    = reg2hw.status_2036.re;


  assign rcache_line[7][245].tag_reg.tag      = reg2hw.tag_2037.q;
  assign rcache_line[7][245].tag_reg.qe       = reg2hw.tag_2037.qe;
  assign rcache_line[7][245].tag_reg.re       = reg2hw.tag_2037.re;
  assign rcache_line[7][245].status_reg.status = reg2hw.status_2037.q;//status_reg_t'(reg2hw.status_2037.q);
  assign rcache_line[7][245].status_reg.qe    = reg2hw.status_2037.qe;
  assign rcache_line[7][245].status_reg.re    = reg2hw.status_2037.re;


  assign rcache_line[7][246].tag_reg.tag      = reg2hw.tag_2038.q;
  assign rcache_line[7][246].tag_reg.qe       = reg2hw.tag_2038.qe;
  assign rcache_line[7][246].tag_reg.re       = reg2hw.tag_2038.re;
  assign rcache_line[7][246].status_reg.status = reg2hw.status_2038.q;//status_reg_t'(reg2hw.status_2038.q);
  assign rcache_line[7][246].status_reg.qe    = reg2hw.status_2038.qe;
  assign rcache_line[7][246].status_reg.re    = reg2hw.status_2038.re;


  assign rcache_line[7][247].tag_reg.tag      = reg2hw.tag_2039.q;
  assign rcache_line[7][247].tag_reg.qe       = reg2hw.tag_2039.qe;
  assign rcache_line[7][247].tag_reg.re       = reg2hw.tag_2039.re;
  assign rcache_line[7][247].status_reg.status = reg2hw.status_2039.q;//status_reg_t'(reg2hw.status_2039.q);
  assign rcache_line[7][247].status_reg.qe    = reg2hw.status_2039.qe;
  assign rcache_line[7][247].status_reg.re    = reg2hw.status_2039.re;


  assign rcache_line[7][248].tag_reg.tag      = reg2hw.tag_2040.q;
  assign rcache_line[7][248].tag_reg.qe       = reg2hw.tag_2040.qe;
  assign rcache_line[7][248].tag_reg.re       = reg2hw.tag_2040.re;
  assign rcache_line[7][248].status_reg.status = reg2hw.status_2040.q;//status_reg_t'(reg2hw.status_2040.q);
  assign rcache_line[7][248].status_reg.qe    = reg2hw.status_2040.qe;
  assign rcache_line[7][248].status_reg.re    = reg2hw.status_2040.re;


  assign rcache_line[7][249].tag_reg.tag      = reg2hw.tag_2041.q;
  assign rcache_line[7][249].tag_reg.qe       = reg2hw.tag_2041.qe;
  assign rcache_line[7][249].tag_reg.re       = reg2hw.tag_2041.re;
  assign rcache_line[7][249].status_reg.status = reg2hw.status_2041.q;//status_reg_t'(reg2hw.status_2041.q);
  assign rcache_line[7][249].status_reg.qe    = reg2hw.status_2041.qe;
  assign rcache_line[7][249].status_reg.re    = reg2hw.status_2041.re;


  assign rcache_line[7][250].tag_reg.tag      = reg2hw.tag_2042.q;
  assign rcache_line[7][250].tag_reg.qe       = reg2hw.tag_2042.qe;
  assign rcache_line[7][250].tag_reg.re       = reg2hw.tag_2042.re;
  assign rcache_line[7][250].status_reg.status = reg2hw.status_2042.q;//status_reg_t'(reg2hw.status_2042.q);
  assign rcache_line[7][250].status_reg.qe    = reg2hw.status_2042.qe;
  assign rcache_line[7][250].status_reg.re    = reg2hw.status_2042.re;


  assign rcache_line[7][251].tag_reg.tag      = reg2hw.tag_2043.q;
  assign rcache_line[7][251].tag_reg.qe       = reg2hw.tag_2043.qe;
  assign rcache_line[7][251].tag_reg.re       = reg2hw.tag_2043.re;
  assign rcache_line[7][251].status_reg.status = reg2hw.status_2043.q;//status_reg_t'(reg2hw.status_2043.q);
  assign rcache_line[7][251].status_reg.qe    = reg2hw.status_2043.qe;
  assign rcache_line[7][251].status_reg.re    = reg2hw.status_2043.re;


  assign rcache_line[7][252].tag_reg.tag      = reg2hw.tag_2044.q;
  assign rcache_line[7][252].tag_reg.qe       = reg2hw.tag_2044.qe;
  assign rcache_line[7][252].tag_reg.re       = reg2hw.tag_2044.re;
  assign rcache_line[7][252].status_reg.status = reg2hw.status_2044.q;//status_reg_t'(reg2hw.status_2044.q);
  assign rcache_line[7][252].status_reg.qe    = reg2hw.status_2044.qe;
  assign rcache_line[7][252].status_reg.re    = reg2hw.status_2044.re;


  assign rcache_line[7][253].tag_reg.tag      = reg2hw.tag_2045.q;
  assign rcache_line[7][253].tag_reg.qe       = reg2hw.tag_2045.qe;
  assign rcache_line[7][253].tag_reg.re       = reg2hw.tag_2045.re;
  assign rcache_line[7][253].status_reg.status = reg2hw.status_2045.q;//status_reg_t'(reg2hw.status_2045.q);
  assign rcache_line[7][253].status_reg.qe    = reg2hw.status_2045.qe;
  assign rcache_line[7][253].status_reg.re    = reg2hw.status_2045.re;


  assign rcache_line[7][254].tag_reg.tag      = reg2hw.tag_2046.q;
  assign rcache_line[7][254].tag_reg.qe       = reg2hw.tag_2046.qe;
  assign rcache_line[7][254].tag_reg.re       = reg2hw.tag_2046.re;
  assign rcache_line[7][254].status_reg.status = reg2hw.status_2046.q;//status_reg_t'(reg2hw.status_2046.q);
  assign rcache_line[7][254].status_reg.qe    = reg2hw.status_2046.qe;
  assign rcache_line[7][254].status_reg.re    = reg2hw.status_2046.re;


  assign rcache_line[7][255].tag_reg.tag      = reg2hw.tag_2047.q;
  assign rcache_line[7][255].tag_reg.qe       = reg2hw.tag_2047.qe;
  assign rcache_line[7][255].tag_reg.re       = reg2hw.tag_2047.re;
  assign rcache_line[7][255].status_reg.status = reg2hw.status_2047.q;//status_reg_t'(reg2hw.status_2047.q);
  assign rcache_line[7][255].status_reg.qe    = reg2hw.status_2047.qe;
  assign rcache_line[7][255].status_reg.re    = reg2hw.status_2047.re;


  logic [NWays-1:0][NSets-1:0] tag_qe; // Valid bits for the tag registers
  logic [NWays-1:0][NSets-1:0] status_qe; // Valid bits for the status registers
  logic [NWays-1:0][NSets-1:0] tag_re; // Valid bits for the tag registers
  logic [NWays-1:0][NSets-1:0] status_re; // Valid bits for the status registers


  always_comb begin
    ram_sw_index = '0; // Default value for the software index
    ram_sw_wdata = '0; // Default value for the software write data
    // Initialize the tag and status valid bits
    for (int i = 0; i < NWays; i++) begin
      for (int j = 0; j < NSets; j++) begin
        if (rcache_line[i][j].tag_reg.qe == 1'b1 && rcache_line[i][j].status_reg.qe == 1'b1) begin
          ram_sw_index = logic'(j);
          ram_sw_wdata = {rcache_line[i][j].status_reg.status, rcache_line[i][j].tag_reg.tag};
        end
      end
    end
  end
  generate
    for (genvar i = 0; i < NWays; i++) begin : gen_way
      assign ram_sw_we[i] = |status_qe[i] & |tag_qe[i]; // Write enable for the tag store
      assign ram_sw_req[i] = (|status_qe[i] & |tag_qe[i]) | (|status_re[i] & |tag_re[i]);
      for (genvar j = 0; j < NSets; j++) begin : gen_set
        assign tag_qe[i][j] = rcache_line[i][j].tag_reg.qe;
        assign status_qe[i][j] = rcache_line[i][j].status_reg.qe;
        assign tag_re[i][j] = rcache_line[i][j].tag_reg.re;
        assign status_re[i][j] = rcache_line[i][j].status_reg.re;
      end

    end
  endgenerate
  // Mux write requests with HW interface
  // ------------------------------------
  assign ram_hw_req = |ram_req_i; // HW request for the way i
  generate
  for (genvar i = 0; i < NWays; i++) begin : gen_mux
      assign ram_req[i] = ram_sw_req[i] || ram_req_i[i]; // Combine SW and HW requests
      assign ram_we[i]  = ram_req_i[i] ? ram_we_i[i] : ram_sw_we[i];
  end
  endgenerate
  // Write and read data
  assign ram_index = ram_hw_req ? ram_addr_i  : ram_sw_index; // Assuming ram_index is the index part of the address
  assign ram_wdata = ram_hw_req ? ram_wdata_i : ram_sw_wdata;
  assign ram_rdata_o = ram_rdata; // Read data from the tag store (no data gating)


  // Read port of memory
  // -------------------
  // Mem has a single read port, so we have that whatever set has the same d.
  // Should not be a problem as d = qs and the correct set output should be selected

  assign hw2reg.tag_0.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_0.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_1.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_2.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_3.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_3.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_4.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_4.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_5.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_5.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_6.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_6.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_7.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_7.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_8.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_8.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_9.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_9.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_10.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_10.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_11.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_11.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_12.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_12.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_13.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_13.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_14.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_14.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_15.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_15.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_16.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_16.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_17.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_17.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_18.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_18.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_19.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_19.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_20.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_20.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_21.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_21.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_22.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_22.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_23.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_23.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_24.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_24.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_25.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_25.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_26.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_26.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_27.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_27.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_28.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_28.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_29.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_29.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_30.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_30.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_31.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_31.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_32.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_32.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_33.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_33.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_34.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_34.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_35.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_35.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_36.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_36.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_37.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_37.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_38.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_38.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_39.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_39.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_40.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_40.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_41.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_41.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_42.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_42.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_43.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_43.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_44.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_44.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_45.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_45.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_46.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_46.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_47.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_47.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_48.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_48.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_49.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_49.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_50.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_50.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_51.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_51.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_52.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_52.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_53.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_53.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_54.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_54.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_55.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_55.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_56.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_56.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_57.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_57.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_58.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_58.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_59.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_59.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_60.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_60.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_61.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_61.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_62.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_62.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_63.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_63.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_64.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_64.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_65.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_65.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_66.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_66.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_67.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_67.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_68.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_68.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_69.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_69.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_70.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_70.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_71.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_71.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_72.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_72.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_73.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_73.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_74.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_74.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_75.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_75.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_76.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_76.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_77.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_77.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_78.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_78.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_79.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_79.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_80.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_80.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_81.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_81.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_82.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_82.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_83.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_83.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_84.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_84.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_85.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_85.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_86.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_86.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_87.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_87.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_88.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_88.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_89.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_89.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_90.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_90.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_91.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_91.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_92.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_92.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_93.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_93.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_94.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_94.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_95.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_95.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_96.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_96.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_97.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_97.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_98.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_98.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_99.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_99.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_100.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_100.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_101.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_101.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_102.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_102.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_103.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_103.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_104.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_104.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_105.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_105.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_106.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_106.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_107.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_107.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_108.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_108.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_109.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_109.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_110.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_110.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_111.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_111.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_112.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_112.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_113.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_113.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_114.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_114.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_115.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_115.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_116.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_116.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_117.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_117.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_118.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_118.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_119.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_119.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_120.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_120.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_121.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_121.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_122.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_122.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_123.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_123.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_124.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_124.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_125.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_125.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_126.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_126.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_127.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_127.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_128.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_128.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_129.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_129.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_130.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_130.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_131.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_131.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_132.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_132.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_133.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_133.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_134.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_134.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_135.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_135.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_136.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_136.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_137.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_137.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_138.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_138.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_139.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_139.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_140.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_140.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_141.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_141.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_142.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_142.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_143.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_143.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_144.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_144.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_145.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_145.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_146.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_146.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_147.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_147.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_148.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_148.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_149.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_149.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_150.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_150.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_151.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_151.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_152.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_152.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_153.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_153.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_154.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_154.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_155.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_155.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_156.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_156.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_157.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_157.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_158.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_158.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_159.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_159.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_160.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_160.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_161.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_161.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_162.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_162.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_163.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_163.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_164.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_164.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_165.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_165.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_166.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_166.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_167.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_167.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_168.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_168.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_169.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_169.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_170.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_170.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_171.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_171.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_172.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_172.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_173.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_173.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_174.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_174.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_175.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_175.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_176.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_176.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_177.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_177.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_178.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_178.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_179.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_179.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_180.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_180.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_181.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_181.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_182.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_182.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_183.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_183.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_184.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_184.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_185.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_185.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_186.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_186.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_187.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_187.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_188.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_188.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_189.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_189.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_190.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_190.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_191.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_191.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_192.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_192.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_193.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_193.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_194.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_194.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_195.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_195.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_196.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_196.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_197.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_197.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_198.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_198.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_199.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_199.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_200.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_200.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_201.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_201.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_202.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_202.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_203.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_203.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_204.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_204.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_205.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_205.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_206.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_206.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_207.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_207.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_208.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_208.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_209.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_209.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_210.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_210.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_211.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_211.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_212.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_212.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_213.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_213.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_214.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_214.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_215.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_215.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_216.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_216.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_217.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_217.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_218.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_218.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_219.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_219.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_220.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_220.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_221.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_221.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_222.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_222.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_223.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_223.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_224.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_224.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_225.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_225.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_226.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_226.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_227.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_227.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_228.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_228.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_229.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_229.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_230.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_230.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_231.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_231.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_232.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_232.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_233.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_233.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_234.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_234.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_235.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_235.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_236.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_236.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_237.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_237.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_238.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_238.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_239.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_239.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_240.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_240.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_241.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_241.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_242.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_242.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_243.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_243.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_244.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_244.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_245.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_245.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_246.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_246.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_247.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_247.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_248.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_248.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_249.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_249.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_250.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_250.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_251.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_251.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_252.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_252.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_253.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_253.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_254.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_254.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_255.d       = ram_rdata[0][DataWidth-1-3:0];
  assign hw2reg.status_255.d    = ram_rdata[0][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_256.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_256.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_257.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_257.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_258.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_258.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_259.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_259.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_260.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_260.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_261.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_261.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_262.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_262.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_263.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_263.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_264.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_264.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_265.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_265.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_266.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_266.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_267.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_267.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_268.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_268.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_269.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_269.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_270.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_270.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_271.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_271.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_272.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_272.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_273.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_273.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_274.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_274.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_275.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_275.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_276.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_276.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_277.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_277.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_278.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_278.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_279.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_279.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_280.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_280.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_281.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_281.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_282.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_282.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_283.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_283.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_284.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_284.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_285.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_285.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_286.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_286.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_287.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_287.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_288.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_288.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_289.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_289.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_290.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_290.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_291.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_291.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_292.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_292.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_293.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_293.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_294.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_294.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_295.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_295.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_296.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_296.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_297.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_297.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_298.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_298.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_299.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_299.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_300.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_300.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_301.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_301.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_302.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_302.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_303.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_303.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_304.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_304.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_305.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_305.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_306.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_306.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_307.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_307.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_308.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_308.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_309.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_309.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_310.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_310.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_311.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_311.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_312.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_312.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_313.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_313.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_314.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_314.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_315.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_315.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_316.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_316.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_317.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_317.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_318.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_318.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_319.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_319.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_320.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_320.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_321.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_321.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_322.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_322.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_323.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_323.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_324.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_324.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_325.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_325.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_326.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_326.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_327.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_327.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_328.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_328.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_329.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_329.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_330.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_330.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_331.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_331.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_332.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_332.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_333.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_333.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_334.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_334.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_335.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_335.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_336.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_336.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_337.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_337.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_338.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_338.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_339.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_339.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_340.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_340.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_341.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_341.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_342.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_342.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_343.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_343.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_344.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_344.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_345.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_345.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_346.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_346.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_347.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_347.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_348.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_348.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_349.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_349.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_350.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_350.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_351.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_351.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_352.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_352.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_353.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_353.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_354.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_354.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_355.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_355.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_356.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_356.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_357.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_357.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_358.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_358.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_359.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_359.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_360.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_360.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_361.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_361.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_362.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_362.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_363.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_363.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_364.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_364.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_365.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_365.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_366.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_366.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_367.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_367.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_368.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_368.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_369.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_369.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_370.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_370.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_371.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_371.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_372.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_372.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_373.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_373.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_374.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_374.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_375.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_375.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_376.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_376.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_377.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_377.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_378.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_378.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_379.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_379.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_380.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_380.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_381.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_381.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_382.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_382.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_383.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_383.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_384.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_384.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_385.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_385.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_386.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_386.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_387.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_387.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_388.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_388.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_389.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_389.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_390.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_390.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_391.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_391.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_392.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_392.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_393.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_393.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_394.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_394.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_395.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_395.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_396.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_396.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_397.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_397.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_398.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_398.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_399.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_399.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_400.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_400.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_401.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_401.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_402.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_402.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_403.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_403.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_404.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_404.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_405.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_405.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_406.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_406.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_407.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_407.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_408.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_408.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_409.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_409.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_410.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_410.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_411.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_411.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_412.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_412.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_413.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_413.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_414.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_414.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_415.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_415.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_416.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_416.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_417.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_417.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_418.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_418.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_419.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_419.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_420.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_420.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_421.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_421.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_422.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_422.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_423.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_423.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_424.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_424.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_425.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_425.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_426.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_426.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_427.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_427.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_428.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_428.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_429.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_429.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_430.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_430.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_431.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_431.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_432.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_432.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_433.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_433.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_434.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_434.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_435.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_435.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_436.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_436.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_437.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_437.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_438.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_438.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_439.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_439.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_440.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_440.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_441.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_441.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_442.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_442.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_443.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_443.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_444.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_444.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_445.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_445.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_446.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_446.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_447.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_447.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_448.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_448.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_449.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_449.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_450.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_450.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_451.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_451.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_452.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_452.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_453.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_453.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_454.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_454.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_455.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_455.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_456.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_456.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_457.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_457.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_458.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_458.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_459.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_459.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_460.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_460.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_461.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_461.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_462.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_462.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_463.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_463.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_464.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_464.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_465.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_465.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_466.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_466.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_467.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_467.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_468.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_468.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_469.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_469.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_470.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_470.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_471.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_471.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_472.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_472.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_473.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_473.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_474.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_474.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_475.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_475.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_476.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_476.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_477.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_477.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_478.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_478.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_479.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_479.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_480.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_480.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_481.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_481.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_482.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_482.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_483.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_483.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_484.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_484.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_485.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_485.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_486.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_486.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_487.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_487.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_488.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_488.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_489.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_489.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_490.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_490.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_491.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_491.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_492.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_492.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_493.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_493.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_494.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_494.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_495.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_495.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_496.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_496.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_497.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_497.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_498.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_498.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_499.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_499.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_500.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_500.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_501.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_501.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_502.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_502.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_503.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_503.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_504.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_504.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_505.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_505.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_506.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_506.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_507.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_507.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_508.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_508.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_509.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_509.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_510.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_510.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_511.d       = ram_rdata[1][DataWidth-1-3:0];
  assign hw2reg.status_511.d    = ram_rdata[1][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_512.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_512.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_513.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_513.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_514.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_514.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_515.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_515.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_516.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_516.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_517.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_517.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_518.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_518.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_519.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_519.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_520.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_520.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_521.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_521.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_522.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_522.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_523.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_523.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_524.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_524.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_525.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_525.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_526.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_526.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_527.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_527.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_528.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_528.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_529.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_529.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_530.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_530.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_531.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_531.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_532.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_532.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_533.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_533.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_534.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_534.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_535.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_535.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_536.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_536.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_537.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_537.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_538.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_538.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_539.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_539.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_540.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_540.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_541.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_541.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_542.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_542.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_543.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_543.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_544.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_544.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_545.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_545.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_546.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_546.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_547.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_547.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_548.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_548.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_549.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_549.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_550.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_550.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_551.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_551.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_552.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_552.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_553.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_553.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_554.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_554.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_555.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_555.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_556.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_556.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_557.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_557.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_558.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_558.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_559.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_559.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_560.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_560.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_561.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_561.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_562.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_562.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_563.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_563.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_564.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_564.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_565.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_565.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_566.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_566.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_567.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_567.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_568.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_568.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_569.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_569.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_570.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_570.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_571.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_571.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_572.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_572.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_573.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_573.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_574.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_574.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_575.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_575.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_576.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_576.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_577.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_577.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_578.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_578.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_579.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_579.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_580.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_580.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_581.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_581.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_582.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_582.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_583.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_583.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_584.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_584.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_585.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_585.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_586.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_586.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_587.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_587.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_588.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_588.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_589.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_589.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_590.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_590.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_591.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_591.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_592.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_592.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_593.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_593.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_594.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_594.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_595.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_595.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_596.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_596.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_597.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_597.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_598.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_598.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_599.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_599.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_600.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_600.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_601.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_601.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_602.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_602.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_603.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_603.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_604.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_604.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_605.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_605.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_606.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_606.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_607.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_607.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_608.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_608.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_609.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_609.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_610.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_610.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_611.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_611.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_612.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_612.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_613.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_613.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_614.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_614.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_615.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_615.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_616.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_616.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_617.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_617.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_618.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_618.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_619.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_619.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_620.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_620.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_621.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_621.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_622.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_622.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_623.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_623.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_624.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_624.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_625.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_625.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_626.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_626.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_627.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_627.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_628.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_628.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_629.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_629.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_630.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_630.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_631.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_631.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_632.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_632.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_633.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_633.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_634.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_634.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_635.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_635.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_636.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_636.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_637.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_637.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_638.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_638.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_639.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_639.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_640.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_640.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_641.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_641.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_642.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_642.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_643.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_643.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_644.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_644.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_645.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_645.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_646.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_646.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_647.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_647.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_648.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_648.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_649.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_649.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_650.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_650.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_651.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_651.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_652.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_652.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_653.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_653.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_654.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_654.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_655.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_655.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_656.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_656.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_657.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_657.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_658.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_658.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_659.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_659.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_660.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_660.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_661.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_661.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_662.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_662.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_663.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_663.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_664.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_664.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_665.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_665.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_666.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_666.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_667.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_667.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_668.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_668.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_669.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_669.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_670.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_670.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_671.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_671.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_672.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_672.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_673.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_673.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_674.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_674.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_675.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_675.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_676.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_676.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_677.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_677.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_678.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_678.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_679.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_679.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_680.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_680.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_681.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_681.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_682.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_682.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_683.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_683.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_684.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_684.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_685.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_685.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_686.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_686.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_687.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_687.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_688.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_688.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_689.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_689.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_690.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_690.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_691.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_691.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_692.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_692.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_693.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_693.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_694.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_694.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_695.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_695.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_696.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_696.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_697.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_697.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_698.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_698.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_699.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_699.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_700.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_700.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_701.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_701.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_702.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_702.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_703.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_703.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_704.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_704.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_705.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_705.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_706.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_706.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_707.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_707.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_708.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_708.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_709.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_709.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_710.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_710.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_711.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_711.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_712.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_712.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_713.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_713.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_714.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_714.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_715.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_715.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_716.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_716.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_717.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_717.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_718.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_718.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_719.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_719.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_720.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_720.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_721.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_721.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_722.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_722.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_723.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_723.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_724.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_724.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_725.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_725.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_726.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_726.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_727.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_727.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_728.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_728.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_729.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_729.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_730.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_730.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_731.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_731.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_732.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_732.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_733.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_733.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_734.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_734.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_735.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_735.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_736.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_736.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_737.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_737.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_738.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_738.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_739.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_739.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_740.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_740.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_741.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_741.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_742.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_742.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_743.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_743.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_744.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_744.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_745.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_745.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_746.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_746.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_747.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_747.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_748.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_748.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_749.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_749.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_750.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_750.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_751.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_751.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_752.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_752.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_753.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_753.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_754.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_754.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_755.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_755.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_756.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_756.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_757.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_757.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_758.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_758.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_759.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_759.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_760.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_760.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_761.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_761.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_762.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_762.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_763.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_763.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_764.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_764.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_765.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_765.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_766.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_766.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_767.d       = ram_rdata[2][DataWidth-1-3:0];
  assign hw2reg.status_767.d    = ram_rdata[2][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_768.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_768.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_769.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_769.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_770.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_770.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_771.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_771.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_772.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_772.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_773.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_773.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_774.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_774.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_775.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_775.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_776.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_776.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_777.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_777.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_778.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_778.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_779.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_779.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_780.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_780.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_781.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_781.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_782.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_782.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_783.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_783.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_784.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_784.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_785.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_785.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_786.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_786.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_787.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_787.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_788.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_788.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_789.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_789.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_790.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_790.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_791.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_791.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_792.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_792.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_793.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_793.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_794.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_794.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_795.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_795.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_796.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_796.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_797.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_797.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_798.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_798.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_799.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_799.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_800.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_800.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_801.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_801.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_802.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_802.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_803.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_803.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_804.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_804.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_805.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_805.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_806.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_806.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_807.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_807.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_808.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_808.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_809.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_809.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_810.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_810.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_811.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_811.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_812.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_812.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_813.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_813.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_814.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_814.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_815.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_815.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_816.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_816.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_817.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_817.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_818.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_818.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_819.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_819.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_820.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_820.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_821.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_821.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_822.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_822.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_823.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_823.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_824.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_824.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_825.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_825.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_826.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_826.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_827.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_827.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_828.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_828.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_829.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_829.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_830.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_830.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_831.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_831.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_832.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_832.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_833.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_833.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_834.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_834.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_835.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_835.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_836.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_836.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_837.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_837.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_838.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_838.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_839.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_839.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_840.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_840.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_841.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_841.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_842.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_842.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_843.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_843.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_844.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_844.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_845.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_845.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_846.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_846.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_847.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_847.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_848.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_848.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_849.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_849.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_850.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_850.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_851.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_851.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_852.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_852.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_853.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_853.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_854.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_854.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_855.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_855.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_856.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_856.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_857.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_857.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_858.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_858.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_859.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_859.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_860.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_860.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_861.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_861.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_862.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_862.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_863.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_863.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_864.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_864.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_865.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_865.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_866.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_866.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_867.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_867.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_868.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_868.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_869.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_869.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_870.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_870.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_871.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_871.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_872.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_872.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_873.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_873.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_874.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_874.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_875.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_875.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_876.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_876.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_877.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_877.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_878.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_878.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_879.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_879.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_880.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_880.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_881.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_881.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_882.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_882.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_883.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_883.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_884.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_884.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_885.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_885.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_886.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_886.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_887.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_887.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_888.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_888.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_889.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_889.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_890.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_890.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_891.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_891.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_892.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_892.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_893.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_893.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_894.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_894.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_895.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_895.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_896.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_896.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_897.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_897.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_898.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_898.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_899.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_899.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_900.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_900.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_901.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_901.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_902.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_902.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_903.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_903.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_904.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_904.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_905.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_905.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_906.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_906.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_907.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_907.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_908.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_908.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_909.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_909.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_910.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_910.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_911.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_911.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_912.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_912.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_913.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_913.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_914.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_914.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_915.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_915.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_916.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_916.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_917.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_917.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_918.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_918.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_919.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_919.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_920.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_920.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_921.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_921.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_922.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_922.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_923.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_923.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_924.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_924.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_925.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_925.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_926.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_926.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_927.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_927.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_928.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_928.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_929.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_929.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_930.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_930.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_931.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_931.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_932.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_932.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_933.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_933.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_934.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_934.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_935.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_935.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_936.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_936.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_937.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_937.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_938.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_938.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_939.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_939.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_940.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_940.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_941.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_941.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_942.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_942.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_943.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_943.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_944.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_944.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_945.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_945.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_946.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_946.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_947.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_947.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_948.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_948.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_949.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_949.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_950.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_950.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_951.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_951.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_952.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_952.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_953.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_953.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_954.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_954.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_955.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_955.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_956.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_956.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_957.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_957.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_958.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_958.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_959.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_959.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_960.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_960.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_961.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_961.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_962.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_962.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_963.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_963.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_964.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_964.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_965.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_965.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_966.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_966.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_967.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_967.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_968.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_968.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_969.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_969.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_970.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_970.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_971.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_971.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_972.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_972.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_973.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_973.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_974.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_974.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_975.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_975.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_976.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_976.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_977.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_977.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_978.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_978.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_979.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_979.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_980.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_980.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_981.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_981.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_982.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_982.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_983.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_983.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_984.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_984.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_985.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_985.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_986.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_986.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_987.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_987.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_988.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_988.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_989.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_989.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_990.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_990.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_991.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_991.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_992.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_992.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_993.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_993.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_994.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_994.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_995.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_995.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_996.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_996.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_997.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_997.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_998.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_998.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_999.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_999.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1000.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1000.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1001.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1001.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1002.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1002.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1003.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1003.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1004.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1004.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1005.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1005.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1006.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1006.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1007.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1007.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1008.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1008.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1009.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1009.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1010.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1010.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1011.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1011.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1012.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1012.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1013.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1013.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1014.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1014.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1015.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1015.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1016.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1016.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1017.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1017.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1018.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1018.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1019.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1019.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1020.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1020.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1021.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1021.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1022.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1022.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1023.d       = ram_rdata[3][DataWidth-1-3:0];
  assign hw2reg.status_1023.d    = ram_rdata[3][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1024.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1024.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1025.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1025.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1026.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1026.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1027.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1027.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1028.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1028.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1029.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1029.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1030.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1030.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1031.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1031.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1032.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1032.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1033.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1033.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1034.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1034.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1035.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1035.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1036.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1036.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1037.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1037.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1038.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1038.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1039.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1039.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1040.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1040.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1041.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1041.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1042.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1042.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1043.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1043.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1044.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1044.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1045.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1045.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1046.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1046.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1047.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1047.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1048.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1048.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1049.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1049.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1050.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1050.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1051.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1051.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1052.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1052.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1053.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1053.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1054.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1054.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1055.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1055.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1056.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1056.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1057.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1057.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1058.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1058.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1059.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1059.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1060.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1060.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1061.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1061.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1062.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1062.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1063.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1063.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1064.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1064.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1065.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1065.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1066.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1066.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1067.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1067.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1068.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1068.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1069.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1069.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1070.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1070.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1071.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1071.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1072.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1072.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1073.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1073.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1074.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1074.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1075.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1075.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1076.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1076.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1077.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1077.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1078.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1078.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1079.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1079.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1080.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1080.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1081.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1081.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1082.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1082.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1083.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1083.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1084.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1084.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1085.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1085.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1086.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1086.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1087.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1087.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1088.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1088.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1089.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1089.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1090.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1090.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1091.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1091.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1092.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1092.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1093.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1093.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1094.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1094.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1095.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1095.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1096.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1096.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1097.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1097.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1098.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1098.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1099.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1099.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1100.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1100.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1101.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1101.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1102.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1102.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1103.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1103.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1104.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1104.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1105.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1105.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1106.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1106.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1107.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1107.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1108.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1108.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1109.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1109.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1110.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1110.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1111.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1111.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1112.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1112.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1113.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1113.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1114.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1114.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1115.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1115.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1116.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1116.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1117.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1117.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1118.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1118.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1119.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1119.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1120.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1120.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1121.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1121.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1122.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1122.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1123.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1123.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1124.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1124.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1125.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1125.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1126.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1126.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1127.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1127.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1128.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1128.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1129.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1129.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1130.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1130.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1131.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1131.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1132.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1132.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1133.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1133.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1134.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1134.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1135.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1135.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1136.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1136.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1137.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1137.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1138.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1138.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1139.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1139.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1140.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1140.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1141.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1141.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1142.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1142.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1143.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1143.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1144.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1144.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1145.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1145.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1146.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1146.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1147.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1147.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1148.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1148.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1149.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1149.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1150.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1150.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1151.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1151.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1152.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1152.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1153.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1153.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1154.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1154.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1155.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1155.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1156.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1156.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1157.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1157.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1158.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1158.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1159.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1159.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1160.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1160.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1161.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1161.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1162.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1162.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1163.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1163.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1164.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1164.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1165.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1165.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1166.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1166.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1167.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1167.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1168.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1168.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1169.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1169.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1170.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1170.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1171.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1171.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1172.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1172.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1173.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1173.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1174.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1174.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1175.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1175.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1176.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1176.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1177.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1177.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1178.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1178.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1179.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1179.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1180.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1180.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1181.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1181.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1182.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1182.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1183.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1183.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1184.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1184.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1185.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1185.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1186.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1186.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1187.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1187.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1188.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1188.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1189.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1189.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1190.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1190.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1191.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1191.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1192.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1192.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1193.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1193.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1194.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1194.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1195.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1195.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1196.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1196.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1197.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1197.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1198.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1198.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1199.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1199.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1200.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1200.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1201.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1201.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1202.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1202.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1203.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1203.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1204.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1204.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1205.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1205.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1206.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1206.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1207.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1207.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1208.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1208.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1209.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1209.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1210.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1210.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1211.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1211.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1212.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1212.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1213.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1213.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1214.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1214.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1215.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1215.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1216.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1216.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1217.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1217.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1218.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1218.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1219.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1219.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1220.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1220.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1221.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1221.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1222.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1222.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1223.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1223.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1224.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1224.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1225.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1225.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1226.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1226.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1227.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1227.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1228.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1228.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1229.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1229.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1230.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1230.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1231.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1231.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1232.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1232.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1233.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1233.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1234.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1234.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1235.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1235.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1236.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1236.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1237.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1237.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1238.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1238.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1239.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1239.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1240.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1240.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1241.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1241.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1242.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1242.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1243.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1243.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1244.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1244.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1245.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1245.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1246.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1246.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1247.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1247.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1248.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1248.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1249.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1249.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1250.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1250.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1251.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1251.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1252.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1252.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1253.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1253.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1254.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1254.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1255.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1255.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1256.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1256.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1257.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1257.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1258.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1258.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1259.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1259.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1260.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1260.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1261.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1261.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1262.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1262.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1263.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1263.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1264.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1264.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1265.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1265.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1266.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1266.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1267.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1267.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1268.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1268.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1269.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1269.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1270.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1270.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1271.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1271.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1272.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1272.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1273.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1273.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1274.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1274.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1275.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1275.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1276.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1276.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1277.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1277.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1278.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1278.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1279.d       = ram_rdata[4][DataWidth-1-3:0];
  assign hw2reg.status_1279.d    = ram_rdata[4][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1280.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1280.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1281.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1281.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1282.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1282.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1283.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1283.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1284.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1284.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1285.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1285.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1286.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1286.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1287.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1287.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1288.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1288.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1289.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1289.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1290.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1290.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1291.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1291.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1292.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1292.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1293.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1293.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1294.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1294.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1295.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1295.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1296.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1296.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1297.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1297.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1298.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1298.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1299.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1299.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1300.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1300.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1301.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1301.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1302.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1302.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1303.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1303.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1304.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1304.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1305.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1305.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1306.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1306.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1307.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1307.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1308.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1308.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1309.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1309.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1310.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1310.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1311.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1311.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1312.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1312.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1313.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1313.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1314.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1314.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1315.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1315.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1316.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1316.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1317.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1317.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1318.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1318.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1319.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1319.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1320.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1320.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1321.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1321.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1322.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1322.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1323.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1323.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1324.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1324.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1325.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1325.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1326.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1326.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1327.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1327.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1328.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1328.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1329.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1329.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1330.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1330.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1331.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1331.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1332.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1332.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1333.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1333.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1334.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1334.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1335.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1335.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1336.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1336.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1337.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1337.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1338.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1338.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1339.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1339.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1340.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1340.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1341.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1341.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1342.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1342.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1343.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1343.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1344.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1344.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1345.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1345.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1346.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1346.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1347.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1347.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1348.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1348.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1349.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1349.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1350.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1350.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1351.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1351.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1352.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1352.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1353.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1353.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1354.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1354.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1355.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1355.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1356.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1356.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1357.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1357.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1358.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1358.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1359.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1359.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1360.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1360.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1361.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1361.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1362.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1362.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1363.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1363.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1364.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1364.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1365.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1365.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1366.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1366.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1367.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1367.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1368.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1368.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1369.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1369.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1370.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1370.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1371.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1371.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1372.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1372.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1373.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1373.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1374.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1374.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1375.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1375.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1376.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1376.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1377.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1377.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1378.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1378.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1379.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1379.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1380.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1380.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1381.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1381.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1382.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1382.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1383.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1383.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1384.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1384.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1385.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1385.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1386.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1386.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1387.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1387.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1388.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1388.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1389.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1389.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1390.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1390.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1391.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1391.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1392.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1392.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1393.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1393.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1394.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1394.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1395.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1395.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1396.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1396.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1397.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1397.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1398.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1398.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1399.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1399.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1400.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1400.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1401.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1401.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1402.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1402.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1403.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1403.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1404.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1404.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1405.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1405.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1406.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1406.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1407.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1407.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1408.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1408.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1409.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1409.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1410.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1410.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1411.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1411.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1412.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1412.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1413.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1413.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1414.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1414.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1415.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1415.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1416.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1416.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1417.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1417.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1418.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1418.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1419.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1419.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1420.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1420.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1421.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1421.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1422.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1422.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1423.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1423.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1424.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1424.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1425.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1425.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1426.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1426.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1427.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1427.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1428.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1428.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1429.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1429.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1430.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1430.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1431.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1431.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1432.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1432.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1433.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1433.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1434.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1434.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1435.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1435.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1436.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1436.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1437.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1437.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1438.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1438.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1439.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1439.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1440.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1440.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1441.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1441.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1442.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1442.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1443.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1443.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1444.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1444.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1445.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1445.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1446.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1446.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1447.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1447.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1448.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1448.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1449.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1449.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1450.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1450.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1451.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1451.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1452.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1452.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1453.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1453.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1454.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1454.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1455.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1455.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1456.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1456.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1457.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1457.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1458.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1458.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1459.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1459.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1460.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1460.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1461.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1461.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1462.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1462.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1463.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1463.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1464.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1464.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1465.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1465.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1466.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1466.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1467.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1467.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1468.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1468.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1469.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1469.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1470.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1470.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1471.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1471.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1472.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1472.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1473.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1473.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1474.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1474.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1475.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1475.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1476.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1476.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1477.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1477.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1478.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1478.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1479.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1479.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1480.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1480.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1481.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1481.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1482.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1482.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1483.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1483.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1484.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1484.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1485.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1485.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1486.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1486.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1487.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1487.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1488.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1488.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1489.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1489.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1490.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1490.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1491.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1491.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1492.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1492.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1493.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1493.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1494.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1494.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1495.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1495.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1496.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1496.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1497.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1497.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1498.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1498.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1499.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1499.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1500.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1500.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1501.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1501.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1502.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1502.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1503.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1503.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1504.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1504.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1505.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1505.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1506.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1506.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1507.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1507.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1508.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1508.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1509.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1509.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1510.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1510.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1511.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1511.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1512.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1512.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1513.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1513.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1514.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1514.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1515.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1515.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1516.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1516.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1517.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1517.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1518.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1518.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1519.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1519.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1520.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1520.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1521.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1521.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1522.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1522.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1523.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1523.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1524.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1524.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1525.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1525.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1526.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1526.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1527.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1527.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1528.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1528.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1529.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1529.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1530.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1530.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1531.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1531.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1532.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1532.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1533.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1533.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1534.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1534.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1535.d       = ram_rdata[5][DataWidth-1-3:0];
  assign hw2reg.status_1535.d    = ram_rdata[5][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1536.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1536.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1537.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1537.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1538.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1538.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1539.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1539.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1540.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1540.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1541.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1541.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1542.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1542.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1543.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1543.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1544.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1544.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1545.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1545.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1546.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1546.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1547.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1547.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1548.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1548.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1549.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1549.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1550.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1550.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1551.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1551.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1552.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1552.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1553.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1553.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1554.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1554.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1555.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1555.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1556.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1556.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1557.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1557.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1558.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1558.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1559.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1559.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1560.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1560.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1561.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1561.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1562.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1562.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1563.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1563.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1564.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1564.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1565.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1565.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1566.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1566.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1567.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1567.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1568.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1568.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1569.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1569.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1570.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1570.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1571.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1571.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1572.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1572.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1573.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1573.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1574.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1574.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1575.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1575.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1576.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1576.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1577.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1577.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1578.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1578.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1579.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1579.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1580.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1580.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1581.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1581.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1582.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1582.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1583.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1583.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1584.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1584.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1585.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1585.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1586.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1586.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1587.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1587.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1588.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1588.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1589.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1589.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1590.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1590.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1591.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1591.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1592.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1592.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1593.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1593.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1594.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1594.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1595.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1595.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1596.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1596.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1597.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1597.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1598.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1598.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1599.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1599.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1600.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1600.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1601.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1601.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1602.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1602.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1603.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1603.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1604.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1604.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1605.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1605.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1606.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1606.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1607.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1607.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1608.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1608.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1609.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1609.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1610.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1610.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1611.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1611.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1612.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1612.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1613.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1613.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1614.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1614.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1615.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1615.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1616.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1616.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1617.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1617.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1618.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1618.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1619.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1619.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1620.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1620.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1621.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1621.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1622.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1622.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1623.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1623.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1624.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1624.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1625.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1625.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1626.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1626.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1627.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1627.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1628.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1628.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1629.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1629.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1630.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1630.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1631.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1631.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1632.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1632.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1633.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1633.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1634.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1634.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1635.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1635.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1636.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1636.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1637.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1637.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1638.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1638.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1639.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1639.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1640.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1640.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1641.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1641.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1642.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1642.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1643.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1643.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1644.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1644.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1645.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1645.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1646.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1646.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1647.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1647.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1648.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1648.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1649.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1649.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1650.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1650.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1651.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1651.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1652.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1652.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1653.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1653.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1654.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1654.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1655.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1655.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1656.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1656.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1657.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1657.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1658.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1658.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1659.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1659.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1660.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1660.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1661.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1661.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1662.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1662.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1663.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1663.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1664.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1664.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1665.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1665.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1666.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1666.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1667.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1667.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1668.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1668.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1669.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1669.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1670.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1670.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1671.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1671.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1672.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1672.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1673.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1673.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1674.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1674.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1675.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1675.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1676.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1676.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1677.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1677.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1678.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1678.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1679.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1679.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1680.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1680.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1681.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1681.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1682.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1682.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1683.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1683.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1684.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1684.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1685.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1685.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1686.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1686.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1687.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1687.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1688.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1688.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1689.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1689.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1690.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1690.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1691.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1691.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1692.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1692.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1693.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1693.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1694.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1694.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1695.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1695.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1696.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1696.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1697.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1697.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1698.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1698.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1699.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1699.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1700.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1700.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1701.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1701.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1702.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1702.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1703.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1703.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1704.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1704.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1705.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1705.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1706.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1706.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1707.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1707.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1708.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1708.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1709.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1709.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1710.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1710.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1711.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1711.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1712.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1712.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1713.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1713.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1714.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1714.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1715.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1715.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1716.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1716.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1717.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1717.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1718.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1718.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1719.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1719.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1720.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1720.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1721.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1721.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1722.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1722.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1723.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1723.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1724.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1724.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1725.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1725.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1726.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1726.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1727.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1727.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1728.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1728.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1729.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1729.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1730.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1730.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1731.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1731.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1732.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1732.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1733.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1733.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1734.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1734.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1735.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1735.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1736.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1736.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1737.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1737.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1738.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1738.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1739.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1739.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1740.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1740.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1741.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1741.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1742.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1742.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1743.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1743.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1744.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1744.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1745.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1745.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1746.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1746.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1747.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1747.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1748.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1748.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1749.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1749.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1750.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1750.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1751.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1751.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1752.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1752.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1753.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1753.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1754.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1754.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1755.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1755.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1756.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1756.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1757.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1757.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1758.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1758.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1759.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1759.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1760.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1760.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1761.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1761.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1762.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1762.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1763.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1763.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1764.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1764.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1765.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1765.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1766.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1766.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1767.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1767.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1768.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1768.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1769.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1769.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1770.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1770.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1771.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1771.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1772.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1772.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1773.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1773.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1774.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1774.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1775.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1775.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1776.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1776.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1777.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1777.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1778.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1778.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1779.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1779.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1780.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1780.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1781.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1781.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1782.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1782.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1783.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1783.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1784.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1784.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1785.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1785.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1786.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1786.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1787.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1787.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1788.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1788.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1789.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1789.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1790.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1790.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1791.d       = ram_rdata[6][DataWidth-1-3:0];
  assign hw2reg.status_1791.d    = ram_rdata[6][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1792.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1792.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1793.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1793.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1794.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1794.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1795.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1795.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1796.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1796.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1797.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1797.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1798.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1798.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1799.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1799.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1800.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1800.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1801.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1801.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1802.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1802.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1803.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1803.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1804.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1804.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1805.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1805.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1806.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1806.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1807.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1807.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1808.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1808.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1809.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1809.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1810.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1810.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1811.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1811.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1812.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1812.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1813.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1813.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1814.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1814.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1815.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1815.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1816.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1816.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1817.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1817.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1818.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1818.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1819.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1819.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1820.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1820.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1821.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1821.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1822.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1822.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1823.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1823.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1824.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1824.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1825.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1825.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1826.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1826.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1827.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1827.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1828.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1828.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1829.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1829.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1830.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1830.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1831.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1831.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1832.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1832.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1833.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1833.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1834.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1834.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1835.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1835.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1836.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1836.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1837.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1837.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1838.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1838.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1839.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1839.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1840.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1840.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1841.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1841.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1842.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1842.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1843.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1843.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1844.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1844.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1845.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1845.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1846.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1846.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1847.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1847.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1848.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1848.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1849.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1849.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1850.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1850.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1851.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1851.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1852.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1852.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1853.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1853.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1854.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1854.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1855.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1855.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1856.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1856.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1857.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1857.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1858.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1858.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1859.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1859.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1860.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1860.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1861.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1861.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1862.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1862.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1863.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1863.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1864.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1864.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1865.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1865.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1866.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1866.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1867.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1867.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1868.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1868.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1869.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1869.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1870.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1870.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1871.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1871.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1872.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1872.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1873.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1873.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1874.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1874.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1875.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1875.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1876.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1876.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1877.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1877.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1878.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1878.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1879.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1879.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1880.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1880.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1881.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1881.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1882.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1882.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1883.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1883.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1884.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1884.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1885.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1885.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1886.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1886.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1887.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1887.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1888.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1888.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1889.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1889.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1890.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1890.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1891.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1891.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1892.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1892.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1893.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1893.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1894.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1894.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1895.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1895.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1896.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1896.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1897.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1897.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1898.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1898.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1899.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1899.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1900.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1900.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1901.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1901.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1902.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1902.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1903.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1903.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1904.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1904.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1905.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1905.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1906.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1906.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1907.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1907.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1908.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1908.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1909.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1909.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1910.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1910.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1911.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1911.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1912.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1912.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1913.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1913.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1914.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1914.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1915.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1915.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1916.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1916.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1917.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1917.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1918.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1918.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1919.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1919.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1920.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1920.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1921.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1921.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1922.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1922.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1923.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1923.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1924.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1924.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1925.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1925.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1926.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1926.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1927.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1927.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1928.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1928.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1929.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1929.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1930.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1930.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1931.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1931.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1932.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1932.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1933.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1933.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1934.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1934.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1935.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1935.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1936.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1936.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1937.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1937.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1938.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1938.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1939.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1939.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1940.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1940.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1941.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1941.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1942.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1942.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1943.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1943.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1944.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1944.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1945.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1945.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1946.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1946.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1947.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1947.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1948.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1948.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1949.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1949.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1950.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1950.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1951.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1951.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1952.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1952.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1953.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1953.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1954.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1954.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1955.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1955.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1956.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1956.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1957.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1957.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1958.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1958.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1959.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1959.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1960.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1960.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1961.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1961.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1962.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1962.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1963.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1963.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1964.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1964.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1965.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1965.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1966.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1966.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1967.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1967.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1968.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1968.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1969.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1969.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1970.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1970.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1971.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1971.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1972.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1972.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1973.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1973.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1974.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1974.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1975.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1975.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1976.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1976.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1977.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1977.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1978.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1978.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1979.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1979.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1980.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1980.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1981.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1981.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1982.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1982.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1983.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1983.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1984.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1984.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1985.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1985.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1986.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1986.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1987.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1987.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1988.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1988.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1989.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1989.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1990.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1990.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1991.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1991.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1992.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1992.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1993.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1993.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1994.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1994.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1995.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1995.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1996.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1996.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1997.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1997.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1998.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1998.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_1999.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_1999.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2000.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2000.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2001.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2001.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2002.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2002.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2003.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2003.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2004.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2004.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2005.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2005.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2006.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2006.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2007.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2007.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2008.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2008.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2009.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2009.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2010.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2010.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2011.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2011.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2012.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2012.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2013.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2013.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2014.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2014.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2015.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2015.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2016.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2016.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2017.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2017.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2018.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2018.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2019.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2019.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2020.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2020.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2021.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2021.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2022.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2022.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2023.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2023.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2024.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2024.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2025.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2025.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2026.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2026.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2027.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2027.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2028.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2028.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2029.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2029.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2030.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2030.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2031.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2031.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2032.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2032.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2033.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2033.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2034.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2034.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2035.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2035.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2036.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2036.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2037.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2037.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2038.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2038.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2039.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2039.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2040.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2040.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2041.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2041.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2042.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2042.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2043.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2043.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2044.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2044.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2045.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2045.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2046.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2046.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  assign hw2reg.tag_2047.d       = ram_rdata[7][DataWidth-1-3:0];
  assign hw2reg.status_2047.d    = ram_rdata[7][DataWidth-1:DataWidth-1-2];

  //-------------
  // Way Memories
  //-------------
  for (genvar i = 0; unsigned'(i) < NWays; i++) begin : gen_tag_macros
    tc_sram #(
      .NumWords    ( NSets                ),
      .DataWidth   ( DataWidth                   ),
      .ByteWidth   ( ByteWidth                   ),
      .NumPorts    ( 32'd1                        ),
      .Latency     ( axi_llc_pkg::TagMacroLatency ),
      .SimInit     ( "none"                       ),
      .PrintSimCfg ( PrintSimCfg                 )
    ) i_tag_store (
      .clk_i,
      .rst_ni,
      .req_i   ( ram_req[i] ),
      .we_i    ( ram_we[i]  ),
      .addr_i  ( ram_index  ),
      .wdata_i ( ram_wdata  ),
      .be_i    ( ram_we[i]  ),
      .rdata_o ( ram_rdata[i] )
    );
 end


  //-------------------
  // Register interface
  //-------------------
  axi_llc_status_reg_top #(
    .reg_req_t(reg_req_t),
    .reg_rsp_t(reg_rsp_t)
  ) axi_llc_status_reg_top_i (
    .clk_i,
    .rst_ni,
    .reg_req_i,
    .reg_rsp_o,
    .reg2hw,
    .hw2reg,
    .devmode_i(1'b1)
  );

endmodule
